* File: sky130_fd_sc_hs__dfsbp_1.pxi.spice
* Created: Thu Aug 27 20:39:03 2020
* 
x_PM_SKY130_FD_SC_HS__DFSBP_1%D N_D_c_270_n N_D_c_275_n N_D_M1007_g N_D_c_276_n
+ N_D_M1000_g D D N_D_c_272_n N_D_c_273_n N_D_c_278_n
+ PM_SKY130_FD_SC_HS__DFSBP_1%D
x_PM_SKY130_FD_SC_HS__DFSBP_1%CLK N_CLK_c_303_n N_CLK_M1033_g N_CLK_c_304_n
+ N_CLK_M1027_g CLK PM_SKY130_FD_SC_HS__DFSBP_1%CLK
x_PM_SKY130_FD_SC_HS__DFSBP_1%A_398_74# N_A_398_74#_M1017_d N_A_398_74#_M1031_d
+ N_A_398_74#_c_336_n N_A_398_74#_c_355_n N_A_398_74#_c_356_n
+ N_A_398_74#_M1024_g N_A_398_74#_M1022_g N_A_398_74#_M1020_g
+ N_A_398_74#_c_357_n N_A_398_74#_M1019_g N_A_398_74#_c_338_n
+ N_A_398_74#_c_358_n N_A_398_74#_c_339_n N_A_398_74#_c_340_n
+ N_A_398_74#_c_359_n N_A_398_74#_c_360_n N_A_398_74#_c_341_n
+ N_A_398_74#_c_342_n N_A_398_74#_c_343_n N_A_398_74#_c_364_n
+ N_A_398_74#_c_365_n N_A_398_74#_c_366_n N_A_398_74#_c_367_n
+ N_A_398_74#_c_368_n N_A_398_74#_c_369_n N_A_398_74#_c_370_n
+ N_A_398_74#_c_371_n N_A_398_74#_c_393_p N_A_398_74#_c_372_n
+ N_A_398_74#_c_373_n N_A_398_74#_c_344_n N_A_398_74#_c_345_n
+ N_A_398_74#_c_346_n N_A_398_74#_c_347_n N_A_398_74#_c_348_n
+ N_A_398_74#_c_375_n N_A_398_74#_c_349_n N_A_398_74#_c_350_n
+ N_A_398_74#_c_376_n N_A_398_74#_c_351_n N_A_398_74#_c_352_n
+ N_A_398_74#_c_353_n PM_SKY130_FD_SC_HS__DFSBP_1%A_398_74#
x_PM_SKY130_FD_SC_HS__DFSBP_1%A_779_380# N_A_779_380#_M1018_s
+ N_A_779_380#_M1003_d N_A_779_380#_c_638_n N_A_779_380#_M1009_g
+ N_A_779_380#_c_632_n N_A_779_380#_M1011_g N_A_779_380#_c_639_n
+ N_A_779_380#_c_633_n N_A_779_380#_c_634_n N_A_779_380#_c_640_n
+ N_A_779_380#_c_641_n N_A_779_380#_c_642_n N_A_779_380#_c_643_n
+ N_A_779_380#_c_635_n N_A_779_380#_c_636_n N_A_779_380#_c_637_n
+ PM_SKY130_FD_SC_HS__DFSBP_1%A_779_380#
x_PM_SKY130_FD_SC_HS__DFSBP_1%A_596_81# N_A_596_81#_M1008_d N_A_596_81#_M1024_d
+ N_A_596_81#_c_740_n N_A_596_81#_c_741_n N_A_596_81#_M1003_g
+ N_A_596_81#_c_723_n N_A_596_81#_M1018_g N_A_596_81#_c_725_n
+ N_A_596_81#_M1012_g N_A_596_81#_c_726_n N_A_596_81#_M1001_g
+ N_A_596_81#_c_727_n N_A_596_81#_c_728_n N_A_596_81#_c_729_n
+ N_A_596_81#_c_730_n N_A_596_81#_c_731_n N_A_596_81#_c_732_n
+ N_A_596_81#_c_733_n N_A_596_81#_c_734_n N_A_596_81#_c_735_n
+ N_A_596_81#_c_744_n N_A_596_81#_c_736_n N_A_596_81#_c_737_n
+ N_A_596_81#_c_738_n N_A_596_81#_c_739_n PM_SKY130_FD_SC_HS__DFSBP_1%A_596_81#
x_PM_SKY130_FD_SC_HS__DFSBP_1%SET_B N_SET_B_c_896_n N_SET_B_c_897_n
+ N_SET_B_M1029_g N_SET_B_M1028_g N_SET_B_M1025_g N_SET_B_c_887_n
+ N_SET_B_c_888_n N_SET_B_c_899_n N_SET_B_M1005_g N_SET_B_c_889_n
+ N_SET_B_c_890_n N_SET_B_c_891_n N_SET_B_c_892_n SET_B N_SET_B_c_905_n
+ N_SET_B_c_894_n N_SET_B_c_895_n PM_SKY130_FD_SC_HS__DFSBP_1%SET_B
x_PM_SKY130_FD_SC_HS__DFSBP_1%A_225_74# N_A_225_74#_M1033_s N_A_225_74#_M1027_s
+ N_A_225_74#_M1017_g N_A_225_74#_c_1034_n N_A_225_74#_M1031_g
+ N_A_225_74#_c_1046_n N_A_225_74#_c_1035_n N_A_225_74#_c_1047_n
+ N_A_225_74#_c_1048_n N_A_225_74#_M1008_g N_A_225_74#_c_1049_n
+ N_A_225_74#_c_1050_n N_A_225_74#_c_1051_n N_A_225_74#_M1023_g
+ N_A_225_74#_c_1052_n N_A_225_74#_M1013_g N_A_225_74#_c_1037_n
+ N_A_225_74#_c_1038_n N_A_225_74#_M1032_g N_A_225_74#_c_1040_n
+ N_A_225_74#_c_1041_n N_A_225_74#_c_1058_n N_A_225_74#_c_1059_n
+ N_A_225_74#_c_1042_n N_A_225_74#_c_1061_n N_A_225_74#_c_1062_n
+ N_A_225_74#_c_1063_n N_A_225_74#_c_1043_n N_A_225_74#_c_1044_n
+ N_A_225_74#_c_1065_n PM_SKY130_FD_SC_HS__DFSBP_1%A_225_74#
x_PM_SKY130_FD_SC_HS__DFSBP_1%A_1510_48# N_A_1510_48#_M1015_d
+ N_A_1510_48#_M1006_s N_A_1510_48#_M1030_g N_A_1510_48#_c_1222_n
+ N_A_1510_48#_c_1223_n N_A_1510_48#_M1002_g N_A_1510_48#_c_1214_n
+ N_A_1510_48#_c_1215_n N_A_1510_48#_c_1216_n N_A_1510_48#_c_1217_n
+ N_A_1510_48#_c_1224_n N_A_1510_48#_c_1218_n N_A_1510_48#_c_1225_n
+ N_A_1510_48#_c_1226_n N_A_1510_48#_c_1219_n N_A_1510_48#_c_1220_n
+ N_A_1510_48#_c_1221_n PM_SKY130_FD_SC_HS__DFSBP_1%A_1510_48#
x_PM_SKY130_FD_SC_HS__DFSBP_1%A_1355_377# N_A_1355_377#_M1020_d
+ N_A_1355_377#_M1013_d N_A_1355_377#_M1005_d N_A_1355_377#_c_1334_n
+ N_A_1355_377#_M1015_g N_A_1355_377#_c_1335_n N_A_1355_377#_c_1336_n
+ N_A_1355_377#_c_1348_n N_A_1355_377#_M1006_g N_A_1355_377#_c_1337_n
+ N_A_1355_377#_M1014_g N_A_1355_377#_c_1349_n N_A_1355_377#_M1016_g
+ N_A_1355_377#_c_1338_n N_A_1355_377#_c_1339_n N_A_1355_377#_M1026_g
+ N_A_1355_377#_c_1341_n N_A_1355_377#_c_1352_n N_A_1355_377#_M1010_g
+ N_A_1355_377#_c_1342_n N_A_1355_377#_c_1343_n N_A_1355_377#_c_1353_n
+ N_A_1355_377#_c_1366_n N_A_1355_377#_c_1354_n N_A_1355_377#_c_1355_n
+ N_A_1355_377#_c_1344_n N_A_1355_377#_c_1356_n N_A_1355_377#_c_1357_n
+ N_A_1355_377#_c_1358_n N_A_1355_377#_c_1359_n N_A_1355_377#_c_1345_n
+ N_A_1355_377#_c_1360_n N_A_1355_377#_c_1346_n N_A_1355_377#_c_1361_n
+ N_A_1355_377#_c_1362_n N_A_1355_377#_c_1363_n N_A_1355_377#_c_1364_n
+ PM_SKY130_FD_SC_HS__DFSBP_1%A_1355_377#
x_PM_SKY130_FD_SC_HS__DFSBP_1%A_2113_74# N_A_2113_74#_M1026_s
+ N_A_2113_74#_M1010_s N_A_2113_74#_c_1534_n N_A_2113_74#_M1004_g
+ N_A_2113_74#_c_1535_n N_A_2113_74#_M1021_g N_A_2113_74#_c_1536_n
+ N_A_2113_74#_c_1537_n N_A_2113_74#_c_1538_n N_A_2113_74#_c_1539_n
+ N_A_2113_74#_c_1540_n N_A_2113_74#_c_1560_n
+ PM_SKY130_FD_SC_HS__DFSBP_1%A_2113_74#
x_PM_SKY130_FD_SC_HS__DFSBP_1%A_27_80# N_A_27_80#_M1007_s N_A_27_80#_M1008_s
+ N_A_27_80#_M1000_s N_A_27_80#_M1024_s N_A_27_80#_c_1589_n N_A_27_80#_c_1590_n
+ N_A_27_80#_c_1595_n N_A_27_80#_c_1596_n N_A_27_80#_c_1597_n
+ N_A_27_80#_c_1591_n N_A_27_80#_c_1592_n N_A_27_80#_c_1599_n
+ N_A_27_80#_c_1641_n N_A_27_80#_c_1593_n PM_SKY130_FD_SC_HS__DFSBP_1%A_27_80#
x_PM_SKY130_FD_SC_HS__DFSBP_1%VPWR N_VPWR_M1000_d N_VPWR_M1027_d N_VPWR_M1009_d
+ N_VPWR_M1029_d N_VPWR_M1002_d N_VPWR_M1006_d N_VPWR_M1010_d N_VPWR_c_1658_n
+ N_VPWR_c_1659_n N_VPWR_c_1660_n N_VPWR_c_1661_n N_VPWR_c_1662_n
+ N_VPWR_c_1663_n N_VPWR_c_1664_n N_VPWR_c_1665_n N_VPWR_c_1666_n VPWR
+ N_VPWR_c_1667_n N_VPWR_c_1668_n N_VPWR_c_1669_n N_VPWR_c_1670_n
+ N_VPWR_c_1671_n N_VPWR_c_1672_n N_VPWR_c_1673_n N_VPWR_c_1657_n
+ N_VPWR_c_1675_n N_VPWR_c_1676_n N_VPWR_c_1677_n N_VPWR_c_1678_n
+ N_VPWR_c_1679_n N_VPWR_c_1680_n PM_SKY130_FD_SC_HS__DFSBP_1%VPWR
x_PM_SKY130_FD_SC_HS__DFSBP_1%Q_N N_Q_N_M1014_d N_Q_N_M1016_d N_Q_N_c_1803_n Q_N
+ Q_N Q_N Q_N Q_N N_Q_N_c_1805_n Q_N PM_SKY130_FD_SC_HS__DFSBP_1%Q_N
x_PM_SKY130_FD_SC_HS__DFSBP_1%Q N_Q_M1021_d N_Q_M1004_d N_Q_c_1834_n
+ N_Q_c_1835_n Q Q Q Q N_Q_c_1836_n PM_SKY130_FD_SC_HS__DFSBP_1%Q
x_PM_SKY130_FD_SC_HS__DFSBP_1%VGND N_VGND_M1007_d N_VGND_M1033_d N_VGND_M1011_d
+ N_VGND_M1028_d N_VGND_M1025_d N_VGND_M1014_s N_VGND_M1026_d N_VGND_c_1854_n
+ N_VGND_c_1855_n N_VGND_c_1856_n N_VGND_c_1857_n N_VGND_c_1858_n
+ N_VGND_c_1859_n N_VGND_c_1860_n N_VGND_c_1861_n N_VGND_c_1862_n
+ N_VGND_c_1863_n N_VGND_c_1864_n VGND N_VGND_c_1865_n N_VGND_c_1866_n
+ N_VGND_c_1867_n N_VGND_c_1868_n N_VGND_c_1869_n N_VGND_c_1870_n
+ N_VGND_c_1871_n N_VGND_c_1872_n N_VGND_c_1873_n N_VGND_c_1874_n
+ N_VGND_c_1875_n PM_SKY130_FD_SC_HS__DFSBP_1%VGND
cc_1 VNB N_D_c_270_n 0.0419528f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_2 VNB N_D_M1007_g 0.0274789f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_3 VNB N_D_c_272_n 0.025337f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_4 VNB N_D_c_273_n 0.00250659f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_5 VNB N_CLK_c_303_n 0.0199636f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.205
cc_6 VNB N_CLK_c_304_n 0.0363814f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.375
cc_7 VNB CLK 0.00902946f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_8 VNB N_A_398_74#_c_336_n 0.0171808f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_9 VNB N_A_398_74#_M1022_g 0.0446757f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_10 VNB N_A_398_74#_c_338_n 0.00892931f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_11 VNB N_A_398_74#_c_339_n 0.0169218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_398_74#_c_340_n 0.00361019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_398_74#_c_341_n 0.00319375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_398_74#_c_342_n 0.00240575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_343_n 0.0254493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_344_n 0.00221741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_345_n 0.0018239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_346_n 0.00460376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_347_n 0.00217282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_348_n 0.0117768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_349_n 0.004676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_350_n 0.0311252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_351_n 0.00489304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_352_n 0.0220283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_353_n 0.0177899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_779_380#_c_632_n 0.0184541f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_27 VNB N_A_779_380#_c_633_n 0.0192733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_779_380#_c_634_n 0.011878f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_29 VNB N_A_779_380#_c_635_n 0.0257785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_779_380#_c_636_n 0.0198399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_779_380#_c_637_n 0.0363032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_596_81#_c_723_n 0.00979214f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_33 VNB N_A_596_81#_M1018_g 0.031127f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_34 VNB N_A_596_81#_c_725_n 0.040633f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_35 VNB N_A_596_81#_c_726_n 0.0189964f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_36 VNB N_A_596_81#_c_727_n 0.00681186f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_37 VNB N_A_596_81#_c_728_n 0.00270325f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_38 VNB N_A_596_81#_c_729_n 0.0121552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_596_81#_c_730_n 0.00622085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_596_81#_c_731_n 0.0124404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_596_81#_c_732_n 0.00316404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_596_81#_c_733_n 0.00348619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_596_81#_c_734_n 5.61828e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_596_81#_c_735_n 0.0192499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_596_81#_c_736_n 0.00641571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_596_81#_c_737_n 0.00220131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_596_81#_c_738_n 0.00333015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_596_81#_c_739_n 0.0357028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_SET_B_M1028_g 0.0548813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_SET_B_M1025_g 0.0362239f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_51 VNB N_SET_B_c_887_n 0.0174323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_SET_B_c_888_n 0.00564647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_SET_B_c_889_n 0.00545817f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.855
cc_54 VNB N_SET_B_c_890_n 0.011778f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_55 VNB N_SET_B_c_891_n 0.00183892f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_56 VNB N_SET_B_c_892_n 9.3748e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB SET_B 6.75578e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SET_B_c_894_n 0.0380623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_SET_B_c_895_n 0.00714345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_225_74#_M1017_g 0.0224618f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_61 VNB N_A_225_74#_c_1034_n 0.0129807f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_62 VNB N_A_225_74#_c_1035_n 0.0320241f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_63 VNB N_A_225_74#_M1008_g 0.0273819f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_64 VNB N_A_225_74#_c_1037_n 0.00999791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_225_74#_c_1038_n 6.48463e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_225_74#_M1032_g 0.0551903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_225_74#_c_1040_n 0.0266488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_225_74#_c_1041_n 0.018475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_225_74#_c_1042_n 0.0104758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_225_74#_c_1043_n 0.0030415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_225_74#_c_1044_n 0.0131011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1510_48#_M1030_g 0.0488917f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_73 VNB N_A_1510_48#_c_1214_n 0.0116397f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_74 VNB N_A_1510_48#_c_1215_n 0.0163178f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_75 VNB N_A_1510_48#_c_1216_n 0.00463124f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.855
cc_76 VNB N_A_1510_48#_c_1217_n 0.00509151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1510_48#_c_1218_n 0.00694629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1510_48#_c_1219_n 0.00256065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1510_48#_c_1220_n 3.86133e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1510_48#_c_1221_n 0.015955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1355_377#_c_1334_n 0.0201771f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.75
cc_82 VNB N_A_1355_377#_c_1335_n 0.0170735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1355_377#_c_1336_n 0.00484113f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.175
cc_84 VNB N_A_1355_377#_c_1337_n 0.022227f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.855
cc_85 VNB N_A_1355_377#_c_1338_n 0.0833563f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.295
cc_86 VNB N_A_1355_377#_c_1339_n 0.0829175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1355_377#_M1026_g 0.0357041f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_88 VNB N_A_1355_377#_c_1341_n 0.00297161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1355_377#_c_1342_n 0.0350006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1355_377#_c_1343_n 0.0121211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1355_377#_c_1344_n 0.00561225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1355_377#_c_1345_n 8.84857e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1355_377#_c_1346_n 2.14136e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2113_74#_c_1534_n 0.041421f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_95 VNB N_A_2113_74#_c_1535_n 0.0226346f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_96 VNB N_A_2113_74#_c_1536_n 0.00643367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2113_74#_c_1537_n 0.00270135f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.175
cc_98 VNB N_A_2113_74#_c_1538_n 8.76539e-19 $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.855
cc_99 VNB N_A_2113_74#_c_1539_n 0.00756196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2113_74#_c_1540_n 0.00315728f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.665
cc_101 VNB N_A_27_80#_c_1589_n 0.0147808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_27_80#_c_1590_n 0.0387846f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_103 VNB N_A_27_80#_c_1591_n 0.00707322f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_104 VNB N_A_27_80#_c_1592_n 0.00791533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_27_80#_c_1593_n 0.00383527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VPWR_c_1657_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_Q_N_c_1803_n 0.00815532f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_108 VNB Q_N 7.79382e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_109 VNB N_Q_N_c_1805_n 0.0117591f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_110 VNB N_Q_c_1834_n 0.0229628f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_111 VNB N_Q_c_1835_n 0.00626527f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_112 VNB N_Q_c_1836_n 0.0284403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1854_n 0.00901699f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_114 VNB N_VGND_c_1855_n 0.0221343f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_115 VNB N_VGND_c_1856_n 0.00564229f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_116 VNB N_VGND_c_1857_n 0.0168622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1858_n 0.00853376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1859_n 0.0134931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1860_n 0.0101134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1861_n 0.0584454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1862_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1863_n 0.0209428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1864_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1865_n 0.0176596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1866_n 0.0413222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1867_n 0.048518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1868_n 0.034271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1869_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1870_n 0.676277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1871_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1872_n 0.00481148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1873_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1874_n 0.0235452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1875_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VPB N_D_c_270_n 0.015544f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_136 VPB N_D_c_275_n 0.0293f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.375
cc_137 VPB N_D_c_276_n 0.0315437f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_138 VPB N_D_c_273_n 0.00196261f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_139 VPB N_D_c_278_n 0.0244664f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_140 VPB N_CLK_c_304_n 0.0231054f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.375
cc_141 VPB N_A_398_74#_c_336_n 0.00445887f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.61
cc_142 VPB N_A_398_74#_c_355_n 0.0480306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_398_74#_c_356_n 0.0149276f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_144 VPB N_A_398_74#_c_357_n 0.065741f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_145 VPB N_A_398_74#_c_358_n 0.00385362f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_146 VPB N_A_398_74#_c_359_n 0.0217877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_398_74#_c_360_n 0.00372642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_398_74#_c_341_n 0.00209213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_398_74#_c_342_n 0.00544086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_398_74#_c_343_n 0.0170949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_398_74#_c_364_n 0.00283177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_398_74#_c_365_n 0.00895942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_398_74#_c_366_n 0.00389271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_398_74#_c_367_n 0.0157592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_398_74#_c_368_n 0.00260538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_398_74#_c_369_n 0.00218562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_398_74#_c_370_n 0.0113219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_398_74#_c_371_n 2.69913e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_398_74#_c_372_n 0.00637994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_398_74#_c_373_n 0.001186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_398_74#_c_345_n 0.00188182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_398_74#_c_375_n 9.20603e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_398_74#_c_376_n 0.00136728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_398_74#_c_351_n 0.00508436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_398_74#_c_352_n 0.014639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_779_380#_c_638_n 0.0147727f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.61
cc_167 VPB N_A_779_380#_c_639_n 0.0103536f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_168 VPB N_A_779_380#_c_640_n 0.0287641f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.01
cc_169 VPB N_A_779_380#_c_641_n 0.00923854f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_170 VPB N_A_779_380#_c_642_n 0.0341146f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_171 VPB N_A_779_380#_c_643_n 0.00377944f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_172 VPB N_A_779_380#_c_636_n 0.00636452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_596_81#_c_740_n 0.0242564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_596_81#_c_741_n 0.0205293f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_175 VPB N_A_596_81#_c_725_n 0.0232119f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_176 VPB N_A_596_81#_c_727_n 0.0104002f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_177 VPB N_A_596_81#_c_744_n 0.00450702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_596_81#_c_736_n 0.00877854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_SET_B_c_896_n 0.0131889f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_180 VPB N_SET_B_c_897_n 0.0208913f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.02
cc_181 VPB N_SET_B_M1028_g 0.00278972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_SET_B_c_899_n 0.0199546f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.175
cc_183 VPB N_SET_B_c_889_n 0.0500303f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.855
cc_184 VPB N_SET_B_c_890_n 0.0176752f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_185 VPB N_SET_B_c_891_n 2.44984e-19 $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_186 VPB N_SET_B_c_892_n 0.00209073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB SET_B 0.00142743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_SET_B_c_905_n 0.0402354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_SET_B_c_895_n 0.00347893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_225_74#_c_1034_n 0.0201055f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_191 VPB N_A_225_74#_c_1046_n 0.0774119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_225_74#_c_1047_n 0.0602166f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_193 VPB N_A_225_74#_c_1048_n 0.0125859f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.01
cc_194 VPB N_A_225_74#_c_1049_n 0.00745764f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_195 VPB N_A_225_74#_c_1050_n 0.0131636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_225_74#_c_1051_n 0.0143883f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_197 VPB N_A_225_74#_c_1052_n 0.230696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_225_74#_M1013_g 0.00984299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_225_74#_c_1037_n 0.0352795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_225_74#_c_1038_n 0.00796722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_225_74#_c_1040_n 6.04301e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_225_74#_c_1041_n 0.0109988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_225_74#_c_1058_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_225_74#_c_1059_n 0.0242482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_225_74#_c_1042_n 0.00236347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_225_74#_c_1061_n 0.00592994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_225_74#_c_1062_n 0.00519182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_225_74#_c_1063_n 0.00500969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_225_74#_c_1043_n 5.21083e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_225_74#_c_1065_n 8.57544e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1510_48#_c_1222_n 0.0230824f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_212 VPB N_A_1510_48#_c_1223_n 0.0203804f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_213 VPB N_A_1510_48#_c_1224_n 0.00688734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1510_48#_c_1225_n 3.23859e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1510_48#_c_1226_n 0.00469097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1510_48#_c_1219_n 0.00737273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1510_48#_c_1221_n 0.0304329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1355_377#_c_1336_n 0.0322333f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.175
cc_219 VPB N_A_1355_377#_c_1348_n 0.0692137f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_220 VPB N_A_1355_377#_c_1349_n 0.0188981f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=2.02
cc_221 VPB N_A_1355_377#_c_1339_n 0.00803755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1355_377#_c_1341_n 0.0078348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1355_377#_c_1352_n 0.0161227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1355_377#_c_1353_n 0.0162513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1355_377#_c_1354_n 0.003873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1355_377#_c_1355_n 0.00226886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1355_377#_c_1356_n 0.00604561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1355_377#_c_1357_n 0.00757363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1355_377#_c_1358_n 0.0192277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1355_377#_c_1359_n 0.00300004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1355_377#_c_1360_n 0.0044999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1355_377#_c_1361_n 0.0012099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1355_377#_c_1362_n 0.00456694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1355_377#_c_1363_n 0.00401902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1355_377#_c_1364_n 0.0107701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_2113_74#_c_1534_n 0.029368f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.61
cc_237 VPB N_A_2113_74#_c_1538_n 0.00971433f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_238 VPB N_A_27_80#_c_1590_n 0.0249205f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_239 VPB N_A_27_80#_c_1595_n 0.027524f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_240 VPB N_A_27_80#_c_1596_n 0.0259099f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=2.02
cc_241 VPB N_A_27_80#_c_1597_n 0.0140698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_27_80#_c_1591_n 0.00269752f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_243 VPB N_A_27_80#_c_1599_n 0.0109364f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_244 VPB N_VPWR_c_1658_n 0.0140914f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_245 VPB N_VPWR_c_1659_n 0.00646119f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_246 VPB N_VPWR_c_1660_n 0.00593216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1661_n 0.00940309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1662_n 0.00805291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1663_n 0.0069087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1664_n 0.012096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1665_n 0.0566956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1666_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1667_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1668_n 0.0215753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1669_n 0.0500512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1670_n 0.029515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1671_n 0.0368168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1672_n 0.0325425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1673_n 0.0193106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1657_n 0.135168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1675_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1676_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1677_n 0.00523428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1678_n 0.00450185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1679_n 0.00653547f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1680_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB Q_N 0.0194901f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_268 VPB Q 0.0523285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_Q_c_1836_n 0.00759307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 N_D_c_272_n N_CLK_c_303_n 0.00207613f $X=0.64 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_271 N_D_c_270_n N_CLK_c_304_n 0.00989855f $X=0.61 $Y=1.825 $X2=0 $Y2=0
cc_272 N_D_c_272_n N_A_225_74#_c_1042_n 0.00683134f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_273 N_D_c_273_n N_A_225_74#_c_1042_n 0.0532484f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_274 N_D_c_270_n N_A_225_74#_c_1062_n 0.00335375f $X=0.61 $Y=1.825 $X2=0 $Y2=0
cc_275 N_D_c_273_n N_A_225_74#_c_1062_n 0.0249554f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_276 N_D_M1007_g N_A_225_74#_c_1044_n 0.00630877f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_277 N_D_M1007_g N_A_27_80#_c_1589_n 0.00146243f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_278 N_D_M1007_g N_A_27_80#_c_1590_n 0.00600966f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_279 N_D_c_272_n N_A_27_80#_c_1590_n 0.0309478f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_280 N_D_c_273_n N_A_27_80#_c_1590_n 0.0697394f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_281 N_D_c_275_n N_A_27_80#_c_1595_n 0.00433476f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_282 N_D_c_276_n N_A_27_80#_c_1595_n 0.00634977f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_283 N_D_c_275_n N_A_27_80#_c_1596_n 0.0215679f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_284 N_D_c_273_n N_A_27_80#_c_1596_n 0.0257673f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_285 N_D_c_278_n N_A_27_80#_c_1596_n 0.00145366f $X=0.64 $Y=1.855 $X2=0 $Y2=0
cc_286 N_D_c_276_n N_VPWR_c_1658_n 0.0121276f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_287 N_D_c_276_n N_VPWR_c_1667_n 0.00413917f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_288 N_D_c_276_n N_VPWR_c_1657_n 0.00859049f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_289 N_D_M1007_g N_VGND_c_1854_n 0.0138986f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_290 N_D_c_272_n N_VGND_c_1854_n 0.00175174f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_291 N_D_c_273_n N_VGND_c_1854_n 0.0220022f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_292 N_D_M1007_g N_VGND_c_1865_n 0.00462012f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_293 N_D_M1007_g N_VGND_c_1870_n 0.00450456f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_294 N_CLK_c_303_n N_A_225_74#_M1017_g 0.0131347f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_295 N_CLK_c_304_n N_A_225_74#_M1017_g 0.014451f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_296 CLK N_A_225_74#_M1017_g 0.00486292f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_297 N_CLK_c_304_n N_A_225_74#_c_1034_n 0.052107f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_298 CLK N_A_225_74#_c_1034_n 9.33251e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_299 N_CLK_c_303_n N_A_225_74#_c_1042_n 0.00324692f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_300 N_CLK_c_304_n N_A_225_74#_c_1042_n 0.0065169f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_301 CLK N_A_225_74#_c_1042_n 0.0287772f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_302 N_CLK_c_304_n N_A_225_74#_c_1061_n 0.00313913f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_303 N_CLK_c_304_n N_A_225_74#_c_1063_n 0.00952984f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_304 N_CLK_c_304_n N_A_225_74#_c_1043_n 9.89907e-19 $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_305 CLK N_A_225_74#_c_1043_n 0.0162663f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_306 N_CLK_c_303_n N_A_225_74#_c_1044_n 0.00765617f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_307 N_CLK_c_304_n N_A_225_74#_c_1044_n 0.00114511f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_308 CLK N_A_225_74#_c_1044_n 0.00762435f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_309 N_CLK_c_304_n N_A_225_74#_c_1065_n 0.00477306f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_310 CLK N_A_225_74#_c_1065_n 0.0369589f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_311 N_CLK_c_304_n N_A_27_80#_c_1596_n 0.0161052f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_312 N_CLK_c_304_n N_VPWR_c_1658_n 0.0112858f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_313 N_CLK_c_304_n N_VPWR_c_1659_n 0.0240415f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_314 N_CLK_c_304_n N_VPWR_c_1668_n 0.0048608f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_315 N_CLK_c_304_n N_VPWR_c_1657_n 0.00480464f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_316 N_CLK_c_303_n N_VGND_c_1854_n 0.00303096f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_317 N_CLK_c_303_n N_VGND_c_1855_n 0.00434272f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_318 N_CLK_c_303_n N_VGND_c_1856_n 0.00300619f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_319 CLK N_VGND_c_1856_n 0.0154902f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_320 N_CLK_c_303_n N_VGND_c_1870_n 0.00825157f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_321 N_A_398_74#_c_364_n N_A_779_380#_c_638_n 0.00261463f $X=3.79 $Y=2.905
+ $X2=0 $Y2=0
cc_322 N_A_398_74#_c_365_n N_A_779_380#_c_638_n 0.00762884f $X=4.61 $Y=2.25
+ $X2=0 $Y2=0
cc_323 N_A_398_74#_c_366_n N_A_779_380#_c_638_n 0.0033251f $X=4.695 $Y=2.905
+ $X2=0 $Y2=0
cc_324 N_A_398_74#_c_375_n N_A_779_380#_c_638_n 0.00281873f $X=3.825 $Y=2.25
+ $X2=0 $Y2=0
cc_325 N_A_398_74#_M1022_g N_A_779_380#_c_632_n 0.0419504f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_326 N_A_398_74#_c_365_n N_A_779_380#_c_639_n 0.0127912f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_327 N_A_398_74#_c_343_n N_A_779_380#_c_634_n 5.49495e-19 $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_328 N_A_398_74#_c_355_n N_A_779_380#_c_640_n 0.00197587f $X=3.03 $Y=1.94
+ $X2=0 $Y2=0
cc_329 N_A_398_74#_c_342_n N_A_779_380#_c_640_n 0.0145213f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_330 N_A_398_74#_c_343_n N_A_779_380#_c_640_n 0.00665252f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_331 N_A_398_74#_c_365_n N_A_779_380#_c_640_n 0.00700346f $X=4.61 $Y=2.25
+ $X2=0 $Y2=0
cc_332 N_A_398_74#_c_375_n N_A_779_380#_c_640_n 0.00138473f $X=3.825 $Y=2.25
+ $X2=0 $Y2=0
cc_333 N_A_398_74#_c_342_n N_A_779_380#_c_641_n 0.0117362f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_334 N_A_398_74#_c_365_n N_A_779_380#_c_641_n 0.0424712f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_335 N_A_398_74#_c_393_p N_A_779_380#_c_641_n 0.00122328f $X=5.95 $Y=2.125
+ $X2=0 $Y2=0
cc_336 N_A_398_74#_c_342_n N_A_779_380#_c_642_n 0.00274395f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_337 N_A_398_74#_c_365_n N_A_779_380#_c_643_n 0.0130522f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_338 N_A_398_74#_c_367_n N_A_779_380#_c_643_n 0.0169124f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_339 N_A_398_74#_c_369_n N_A_779_380#_c_643_n 0.0318348f $X=5.455 $Y=2.905
+ $X2=0 $Y2=0
cc_340 N_A_398_74#_c_371_n N_A_779_380#_c_643_n 0.0138639f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_341 N_A_398_74#_c_393_p N_A_779_380#_c_643_n 0.00362126f $X=5.95 $Y=2.125
+ $X2=0 $Y2=0
cc_342 N_A_398_74#_c_342_n N_A_779_380#_c_636_n 0.00137731f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_343 N_A_398_74#_c_343_n N_A_779_380#_c_636_n 0.00875274f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_344 N_A_398_74#_M1022_g N_A_779_380#_c_637_n 0.00279772f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_345 N_A_398_74#_c_339_n N_A_596_81#_M1008_d 2.28826e-19 $X=3.025 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_346 N_A_398_74#_c_348_n N_A_596_81#_M1008_d 0.00589878f $X=3.03 $Y=1.435
+ $X2=-0.19 $Y2=-0.245
cc_347 N_A_398_74#_c_365_n N_A_596_81#_c_741_n 0.0040112f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_348 N_A_398_74#_c_366_n N_A_596_81#_c_741_n 0.0114545f $X=4.695 $Y=2.905
+ $X2=0 $Y2=0
cc_349 N_A_398_74#_c_367_n N_A_596_81#_c_741_n 0.0038873f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_350 N_A_398_74#_c_369_n N_A_596_81#_c_741_n 6.20244e-19 $X=5.455 $Y=2.905
+ $X2=0 $Y2=0
cc_351 N_A_398_74#_c_369_n N_A_596_81#_c_725_n 0.00286832f $X=5.455 $Y=2.905
+ $X2=0 $Y2=0
cc_352 N_A_398_74#_c_370_n N_A_596_81#_c_725_n 0.00575577f $X=5.865 $Y=2.21
+ $X2=0 $Y2=0
cc_353 N_A_398_74#_c_393_p N_A_596_81#_c_725_n 0.00858315f $X=5.95 $Y=2.125
+ $X2=0 $Y2=0
cc_354 N_A_398_74#_c_372_n N_A_596_81#_c_725_n 0.0171084f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_355 N_A_398_74#_c_373_n N_A_596_81#_c_725_n 6.8465e-19 $X=6.035 $Y=1.705
+ $X2=0 $Y2=0
cc_356 N_A_398_74#_c_345_n N_A_596_81#_c_725_n 0.00587485f $X=6.52 $Y=1.62 $X2=0
+ $Y2=0
cc_357 N_A_398_74#_c_349_n N_A_596_81#_c_725_n 0.00226831f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_358 N_A_398_74#_c_350_n N_A_596_81#_c_725_n 0.0174522f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_359 N_A_398_74#_c_344_n N_A_596_81#_c_726_n 0.0078857f $X=6.52 $Y=1.12 $X2=0
+ $Y2=0
cc_360 N_A_398_74#_c_347_n N_A_596_81#_c_726_n 0.00154379f $X=6.605 $Y=0.34
+ $X2=0 $Y2=0
cc_361 N_A_398_74#_c_353_n N_A_596_81#_c_726_n 0.0242288f $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_362 N_A_398_74#_M1022_g N_A_596_81#_c_728_n 0.0102403f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_363 N_A_398_74#_c_339_n N_A_596_81#_c_728_n 0.00340526f $X=3.025 $Y=0.34
+ $X2=0 $Y2=0
cc_364 N_A_398_74#_c_348_n N_A_596_81#_c_728_n 0.0344948f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_365 N_A_398_74#_M1022_g N_A_596_81#_c_729_n 0.0134244f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_366 N_A_398_74#_c_342_n N_A_596_81#_c_729_n 0.012122f $X=3.825 $Y=1.525 $X2=0
+ $Y2=0
cc_367 N_A_398_74#_c_343_n N_A_596_81#_c_729_n 0.00250611f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_368 N_A_398_74#_M1022_g N_A_596_81#_c_730_n 0.00262599f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_369 N_A_398_74#_c_342_n N_A_596_81#_c_730_n 0.00546472f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_370 N_A_398_74#_c_343_n N_A_596_81#_c_730_n 6.63991e-19 $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_371 N_A_398_74#_c_342_n N_A_596_81#_c_732_n 0.0140304f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_372 N_A_398_74#_c_343_n N_A_596_81#_c_732_n 0.00182995f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_373 N_A_398_74#_c_365_n N_A_596_81#_c_732_n 0.00421951f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_374 N_A_398_74#_c_373_n N_A_596_81#_c_735_n 0.00241845f $X=6.035 $Y=1.705
+ $X2=0 $Y2=0
cc_375 N_A_398_74#_c_356_n N_A_596_81#_c_744_n 0.00240648f $X=3.065 $Y=2.24
+ $X2=0 $Y2=0
cc_376 N_A_398_74#_c_359_n N_A_596_81#_c_744_n 0.0238882f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_377 N_A_398_74#_c_341_n N_A_596_81#_c_744_n 0.00142555f $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_378 N_A_398_74#_c_364_n N_A_596_81#_c_744_n 0.0296994f $X=3.79 $Y=2.905 $X2=0
+ $Y2=0
cc_379 N_A_398_74#_c_352_n N_A_596_81#_c_744_n 0.00439492f $X=3.59 $Y=1.525
+ $X2=0 $Y2=0
cc_380 N_A_398_74#_c_355_n N_A_596_81#_c_736_n 0.00933519f $X=3.03 $Y=1.94 $X2=0
+ $Y2=0
cc_381 N_A_398_74#_c_356_n N_A_596_81#_c_736_n 5.4541e-19 $X=3.065 $Y=2.24 $X2=0
+ $Y2=0
cc_382 N_A_398_74#_M1022_g N_A_596_81#_c_736_n 0.00867403f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_383 N_A_398_74#_c_342_n N_A_596_81#_c_736_n 0.0599451f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_384 N_A_398_74#_c_348_n N_A_596_81#_c_736_n 0.0778256f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_385 N_A_398_74#_c_375_n N_A_596_81#_c_736_n 0.0138873f $X=3.825 $Y=2.25 $X2=0
+ $Y2=0
cc_386 N_A_398_74#_c_352_n N_A_596_81#_c_736_n 0.0189266f $X=3.59 $Y=1.525 $X2=0
+ $Y2=0
cc_387 N_A_398_74#_M1022_g N_A_596_81#_c_737_n 0.00408316f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_388 N_A_398_74#_c_348_n N_A_596_81#_c_737_n 0.0143574f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_389 N_A_398_74#_c_352_n N_A_596_81#_c_737_n 0.0018726f $X=3.59 $Y=1.525 $X2=0
+ $Y2=0
cc_390 N_A_398_74#_c_372_n N_A_596_81#_c_738_n 0.014583f $X=6.435 $Y=1.705 $X2=0
+ $Y2=0
cc_391 N_A_398_74#_c_373_n N_A_596_81#_c_738_n 0.00671279f $X=6.035 $Y=1.705
+ $X2=0 $Y2=0
cc_392 N_A_398_74#_c_349_n N_A_596_81#_c_738_n 0.0267149f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_393 N_A_398_74#_c_350_n N_A_596_81#_c_738_n 3.11291e-19 $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_394 N_A_398_74#_c_371_n N_SET_B_c_896_n 0.00295786f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_395 N_A_398_74#_c_393_p N_SET_B_c_896_n 0.00164437f $X=5.95 $Y=2.125 $X2=0
+ $Y2=0
cc_396 N_A_398_74#_c_367_n N_SET_B_c_897_n 0.00146141f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_397 N_A_398_74#_c_369_n N_SET_B_c_897_n 0.0174108f $X=5.455 $Y=2.905 $X2=0
+ $Y2=0
cc_398 N_A_398_74#_c_371_n N_SET_B_c_897_n 0.00554186f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_399 N_A_398_74#_c_373_n N_SET_B_M1028_g 0.00122003f $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_400 N_A_398_74#_c_346_n N_SET_B_M1025_g 4.68011e-19 $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_401 N_A_398_74#_c_351_n N_SET_B_M1025_g 0.00193116f $X=7.395 $Y=2.02 $X2=0
+ $Y2=0
cc_402 N_A_398_74#_c_357_n N_SET_B_c_890_n 2.50329e-19 $X=7.51 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_398_74#_c_370_n N_SET_B_c_890_n 0.00636507f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_404 N_A_398_74#_c_372_n N_SET_B_c_890_n 0.0372227f $X=6.435 $Y=1.705 $X2=0
+ $Y2=0
cc_405 N_A_398_74#_c_373_n N_SET_B_c_890_n 0.0130627f $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_406 N_A_398_74#_c_345_n N_SET_B_c_890_n 0.0035869f $X=6.52 $Y=1.62 $X2=0
+ $Y2=0
cc_407 N_A_398_74#_c_349_n N_SET_B_c_890_n 0.0116123f $X=6.715 $Y=1.285 $X2=0
+ $Y2=0
cc_408 N_A_398_74#_c_350_n N_SET_B_c_890_n 0.00369024f $X=6.715 $Y=1.285 $X2=0
+ $Y2=0
cc_409 N_A_398_74#_c_376_n N_SET_B_c_890_n 0.00592462f $X=7.395 $Y=2.185 $X2=0
+ $Y2=0
cc_410 N_A_398_74#_c_351_n N_SET_B_c_890_n 0.0190815f $X=7.395 $Y=2.02 $X2=0
+ $Y2=0
cc_411 N_A_398_74#_c_370_n N_SET_B_c_891_n 6.26369e-19 $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_412 N_A_398_74#_c_371_n N_SET_B_c_891_n 0.00191865f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_413 N_A_398_74#_c_373_n N_SET_B_c_891_n 3.52044e-19 $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_414 N_A_398_74#_c_370_n N_SET_B_c_892_n 0.0111106f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_415 N_A_398_74#_c_371_n N_SET_B_c_892_n 0.0104469f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_416 N_A_398_74#_c_393_p N_SET_B_c_892_n 0.0120255f $X=5.95 $Y=2.125 $X2=0
+ $Y2=0
cc_417 N_A_398_74#_c_373_n N_SET_B_c_892_n 0.0121378f $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_418 N_A_398_74#_c_370_n N_SET_B_c_905_n 0.00106941f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_419 N_A_398_74#_c_371_n N_SET_B_c_905_n 3.95737e-19 $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_420 N_A_398_74#_c_393_p N_SET_B_c_905_n 0.00134198f $X=5.95 $Y=2.125 $X2=0
+ $Y2=0
cc_421 N_A_398_74#_c_338_n N_A_225_74#_M1017_g 0.00167653f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_422 N_A_398_74#_c_340_n N_A_225_74#_M1017_g 0.00266901f $X=2.295 $Y=0.34
+ $X2=0 $Y2=0
cc_423 N_A_398_74#_c_358_n N_A_225_74#_c_1034_n 0.0048124f $X=2.19 $Y=2.565
+ $X2=0 $Y2=0
cc_424 N_A_398_74#_c_360_n N_A_225_74#_c_1034_n 0.00130182f $X=2.355 $Y=2.99
+ $X2=0 $Y2=0
cc_425 N_A_398_74#_c_355_n N_A_225_74#_c_1046_n 0.0163444f $X=3.03 $Y=1.94 $X2=0
+ $Y2=0
cc_426 N_A_398_74#_c_356_n N_A_225_74#_c_1046_n 0.0111889f $X=3.065 $Y=2.24
+ $X2=0 $Y2=0
cc_427 N_A_398_74#_c_358_n N_A_225_74#_c_1046_n 0.00734636f $X=2.19 $Y=2.565
+ $X2=0 $Y2=0
cc_428 N_A_398_74#_c_359_n N_A_225_74#_c_1046_n 0.0117161f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_429 N_A_398_74#_c_341_n N_A_225_74#_c_1046_n 3.43168e-19 $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_430 N_A_398_74#_c_336_n N_A_225_74#_c_1035_n 0.00655065f $X=3.03 $Y=1.69
+ $X2=0 $Y2=0
cc_431 N_A_398_74#_c_341_n N_A_225_74#_c_1035_n 8.57179e-19 $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_432 N_A_398_74#_c_356_n N_A_225_74#_c_1047_n 0.00882199f $X=3.065 $Y=2.24
+ $X2=0 $Y2=0
cc_433 N_A_398_74#_c_359_n N_A_225_74#_c_1047_n 0.0147556f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_434 N_A_398_74#_M1022_g N_A_225_74#_M1008_g 0.00834991f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_c_338_n N_A_225_74#_M1008_g 0.00333039f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_436 N_A_398_74#_c_339_n N_A_225_74#_M1008_g 0.0158823f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_437 N_A_398_74#_c_348_n N_A_225_74#_M1008_g 0.00854965f $X=3.03 $Y=1.435
+ $X2=0 $Y2=0
cc_438 N_A_398_74#_c_356_n N_A_225_74#_c_1049_n 0.00216849f $X=3.065 $Y=2.24
+ $X2=0 $Y2=0
cc_439 N_A_398_74#_c_364_n N_A_225_74#_c_1049_n 0.00286544f $X=3.79 $Y=2.905
+ $X2=0 $Y2=0
cc_440 N_A_398_74#_c_359_n N_A_225_74#_c_1050_n 0.0175868f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_441 N_A_398_74#_c_355_n N_A_225_74#_c_1051_n 0.00178403f $X=3.03 $Y=1.94
+ $X2=0 $Y2=0
cc_442 N_A_398_74#_c_356_n N_A_225_74#_c_1051_n 0.0107674f $X=3.065 $Y=2.24
+ $X2=0 $Y2=0
cc_443 N_A_398_74#_c_364_n N_A_225_74#_c_1051_n 0.00443587f $X=3.79 $Y=2.905
+ $X2=0 $Y2=0
cc_444 N_A_398_74#_c_375_n N_A_225_74#_c_1051_n 0.00115602f $X=3.825 $Y=2.25
+ $X2=0 $Y2=0
cc_445 N_A_398_74#_c_352_n N_A_225_74#_c_1051_n 0.00476032f $X=3.59 $Y=1.525
+ $X2=0 $Y2=0
cc_446 N_A_398_74#_c_359_n N_A_225_74#_c_1052_n 0.00535373f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_447 N_A_398_74#_c_367_n N_A_225_74#_c_1052_n 0.0130411f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_448 N_A_398_74#_c_368_n N_A_225_74#_c_1052_n 0.00420304f $X=4.78 $Y=2.99
+ $X2=0 $Y2=0
cc_449 N_A_398_74#_c_357_n N_A_225_74#_M1013_g 0.00654176f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_450 N_A_398_74#_c_351_n N_A_225_74#_M1013_g 2.36761e-19 $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_451 N_A_398_74#_c_357_n N_A_225_74#_c_1037_n 0.00534578f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_452 N_A_398_74#_c_376_n N_A_225_74#_c_1037_n 6.10091e-19 $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_372_n N_A_225_74#_c_1038_n 0.00158247f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_454 N_A_398_74#_c_349_n N_A_225_74#_c_1038_n 0.00133533f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_455 N_A_398_74#_c_350_n N_A_225_74#_c_1038_n 0.0194882f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_456 N_A_398_74#_c_345_n N_A_225_74#_M1032_g 7.76595e-19 $X=6.52 $Y=1.62 $X2=0
+ $Y2=0
cc_457 N_A_398_74#_c_346_n N_A_225_74#_M1032_g 0.0120073f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_458 N_A_398_74#_c_349_n N_A_225_74#_M1032_g 3.48236e-19 $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_459 N_A_398_74#_c_350_n N_A_225_74#_M1032_g 0.0149282f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_460 N_A_398_74#_c_351_n N_A_225_74#_M1032_g 0.0115834f $X=7.395 $Y=2.02 $X2=0
+ $Y2=0
cc_461 N_A_398_74#_c_353_n N_A_225_74#_M1032_g 0.0215718f $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_462 N_A_398_74#_c_336_n N_A_225_74#_c_1040_n 0.0130852f $X=3.03 $Y=1.69 $X2=0
+ $Y2=0
cc_463 N_A_398_74#_c_338_n N_A_225_74#_c_1040_n 9.09054e-19 $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_464 N_A_398_74#_c_339_n N_A_225_74#_c_1040_n 0.0034994f $X=3.025 $Y=0.34
+ $X2=0 $Y2=0
cc_465 N_A_398_74#_c_341_n N_A_225_74#_c_1040_n 3.43168e-19 $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_466 N_A_398_74#_c_348_n N_A_225_74#_c_1040_n 7.05733e-19 $X=3.03 $Y=1.435
+ $X2=0 $Y2=0
cc_467 N_A_398_74#_c_338_n N_A_225_74#_c_1041_n 0.00169375f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_357_n N_A_225_74#_c_1059_n 0.00309579f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_469 N_A_398_74#_M1031_d N_A_225_74#_c_1063_n 0.00302182f $X=2.04 $Y=1.79
+ $X2=0 $Y2=0
cc_470 N_A_398_74#_c_338_n N_A_225_74#_c_1043_n 0.0218452f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_471 N_A_398_74#_c_346_n N_A_1510_48#_M1030_g 0.00449224f $X=7.39 $Y=0.34
+ $X2=0 $Y2=0
cc_472 N_A_398_74#_c_351_n N_A_1510_48#_M1030_g 0.0218033f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_473 N_A_398_74#_c_357_n N_A_1510_48#_c_1222_n 0.0215016f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_474 N_A_398_74#_c_376_n N_A_1510_48#_c_1222_n 4.62583e-19 $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_475 N_A_398_74#_c_351_n N_A_1510_48#_c_1222_n 0.00323148f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_476 N_A_398_74#_c_357_n N_A_1510_48#_c_1223_n 0.0285542f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_477 N_A_398_74#_c_351_n N_A_1510_48#_c_1214_n 0.0541231f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_478 N_A_398_74#_c_351_n N_A_1510_48#_c_1216_n 0.0117101f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_479 N_A_398_74#_c_357_n N_A_1510_48#_c_1221_n 0.00165228f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_480 N_A_398_74#_c_351_n N_A_1510_48#_c_1221_n 0.00609625f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_481 N_A_398_74#_c_346_n N_A_1355_377#_M1020_d 0.00260527f $X=7.39 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_482 N_A_398_74#_c_357_n N_A_1355_377#_c_1366_n 0.00530981f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_483 N_A_398_74#_c_376_n N_A_1355_377#_c_1366_n 0.0139926f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_484 N_A_398_74#_c_357_n N_A_1355_377#_c_1354_n 0.00458462f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_485 N_A_398_74#_c_376_n N_A_1355_377#_c_1354_n 0.0260807f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_486 N_A_398_74#_c_372_n N_A_1355_377#_c_1344_n 0.00151891f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_487 N_A_398_74#_c_344_n N_A_1355_377#_c_1344_n 0.0057326f $X=6.52 $Y=1.12
+ $X2=0 $Y2=0
cc_488 N_A_398_74#_c_345_n N_A_1355_377#_c_1344_n 0.00625163f $X=6.52 $Y=1.62
+ $X2=0 $Y2=0
cc_489 N_A_398_74#_c_349_n N_A_1355_377#_c_1344_n 0.025349f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_490 N_A_398_74#_c_350_n N_A_1355_377#_c_1344_n 0.00103124f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_491 N_A_398_74#_c_351_n N_A_1355_377#_c_1344_n 0.0536421f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_492 N_A_398_74#_c_353_n N_A_1355_377#_c_1344_n 0.00145074f $X=6.715 $Y=1.12
+ $X2=0 $Y2=0
cc_493 N_A_398_74#_c_357_n N_A_1355_377#_c_1360_n 5.39738e-19 $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_494 N_A_398_74#_c_372_n N_A_1355_377#_c_1360_n 0.00643961f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_495 N_A_398_74#_c_349_n N_A_1355_377#_c_1360_n 0.00247197f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_496 N_A_398_74#_c_350_n N_A_1355_377#_c_1360_n 2.07025e-19 $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_497 N_A_398_74#_c_376_n N_A_1355_377#_c_1360_n 0.00406811f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_498 N_A_398_74#_c_351_n N_A_1355_377#_c_1360_n 0.0199168f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_499 N_A_398_74#_c_346_n N_A_1355_377#_c_1346_n 0.0232966f $X=7.39 $Y=0.34
+ $X2=0 $Y2=0
cc_500 N_A_398_74#_c_349_n N_A_1355_377#_c_1346_n 0.0051699f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_501 N_A_398_74#_c_350_n N_A_1355_377#_c_1346_n 0.00163857f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_502 N_A_398_74#_c_351_n N_A_1355_377#_c_1346_n 0.0250923f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_503 N_A_398_74#_c_353_n N_A_1355_377#_c_1346_n 0.0040576f $X=6.715 $Y=1.12
+ $X2=0 $Y2=0
cc_504 N_A_398_74#_c_357_n N_A_1355_377#_c_1361_n 0.00697269f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_505 N_A_398_74#_c_357_n N_A_1355_377#_c_1362_n 0.010218f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_506 N_A_398_74#_c_357_n N_A_1355_377#_c_1363_n 0.00670998f $X=7.51 $Y=2.465
+ $X2=0 $Y2=0
cc_507 N_A_398_74#_c_376_n N_A_1355_377#_c_1363_n 0.0218418f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_508 N_A_398_74#_c_339_n N_A_27_80#_M1008_s 0.00233785f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_509 N_A_398_74#_M1031_d N_A_27_80#_c_1597_n 0.00506706f $X=2.04 $Y=1.79 $X2=0
+ $Y2=0
cc_510 N_A_398_74#_c_355_n N_A_27_80#_c_1597_n 0.00322323f $X=3.03 $Y=1.94 $X2=0
+ $Y2=0
cc_511 N_A_398_74#_c_356_n N_A_27_80#_c_1597_n 0.00588528f $X=3.065 $Y=2.24
+ $X2=0 $Y2=0
cc_512 N_A_398_74#_c_358_n N_A_27_80#_c_1597_n 0.0470269f $X=2.19 $Y=2.565 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_359_n N_A_27_80#_c_1597_n 0.0381815f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_c_341_n N_A_27_80#_c_1597_n 0.0147263f $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_c_336_n N_A_27_80#_c_1591_n 0.00427076f $X=3.03 $Y=1.69 $X2=0
+ $Y2=0
cc_516 N_A_398_74#_c_341_n N_A_27_80#_c_1591_n 0.0468227f $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_348_n N_A_27_80#_c_1591_n 0.0274015f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_518 N_A_398_74#_c_338_n N_A_27_80#_c_1593_n 0.0340448f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_c_339_n N_A_27_80#_c_1593_n 0.0199805f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_520 N_A_398_74#_c_348_n N_A_27_80#_c_1593_n 0.0100954f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_521 N_A_398_74#_c_365_n N_VPWR_M1009_d 0.0104455f $X=4.61 $Y=2.25 $X2=0 $Y2=0
cc_522 N_A_398_74#_c_366_n N_VPWR_M1009_d 0.00817577f $X=4.695 $Y=2.905 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_c_369_n N_VPWR_M1029_d 0.00509113f $X=5.455 $Y=2.905 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_370_n N_VPWR_M1029_d 0.00602065f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_393_p N_VPWR_M1029_d 0.00982325f $X=5.95 $Y=2.125 $X2=0
+ $Y2=0
cc_526 N_A_398_74#_c_372_n N_VPWR_M1029_d 8.09396e-19 $X=6.435 $Y=1.705 $X2=0
+ $Y2=0
cc_527 N_A_398_74#_c_373_n N_VPWR_M1029_d 8.27891e-19 $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_528 N_A_398_74#_c_358_n N_VPWR_c_1659_n 0.0251101f $X=2.19 $Y=2.565 $X2=0
+ $Y2=0
cc_529 N_A_398_74#_c_360_n N_VPWR_c_1659_n 0.0128267f $X=2.355 $Y=2.99 $X2=0
+ $Y2=0
cc_530 N_A_398_74#_c_359_n N_VPWR_c_1660_n 0.0152339f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_531 N_A_398_74#_c_364_n N_VPWR_c_1660_n 0.0219178f $X=3.79 $Y=2.905 $X2=0
+ $Y2=0
cc_532 N_A_398_74#_c_365_n N_VPWR_c_1660_n 0.0272218f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_533 N_A_398_74#_c_366_n N_VPWR_c_1660_n 0.0314632f $X=4.695 $Y=2.905 $X2=0
+ $Y2=0
cc_534 N_A_398_74#_c_368_n N_VPWR_c_1660_n 0.0152343f $X=4.78 $Y=2.99 $X2=0
+ $Y2=0
cc_535 N_A_398_74#_c_367_n N_VPWR_c_1661_n 0.0150706f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_536 N_A_398_74#_c_369_n N_VPWR_c_1661_n 0.0340923f $X=5.455 $Y=2.905 $X2=0
+ $Y2=0
cc_537 N_A_398_74#_c_370_n N_VPWR_c_1661_n 0.0280035f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_538 N_A_398_74#_c_372_n N_VPWR_c_1661_n 3.88767e-19 $X=6.435 $Y=1.705 $X2=0
+ $Y2=0
cc_539 N_A_398_74#_c_357_n N_VPWR_c_1665_n 0.00328026f $X=7.51 $Y=2.465 $X2=0
+ $Y2=0
cc_540 N_A_398_74#_c_359_n N_VPWR_c_1669_n 0.0975181f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_541 N_A_398_74#_c_360_n N_VPWR_c_1669_n 0.0179117f $X=2.355 $Y=2.99 $X2=0
+ $Y2=0
cc_542 N_A_398_74#_c_367_n N_VPWR_c_1670_n 0.0495251f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_543 N_A_398_74#_c_368_n N_VPWR_c_1670_n 0.0115893f $X=4.78 $Y=2.99 $X2=0
+ $Y2=0
cc_544 N_A_398_74#_c_357_n N_VPWR_c_1657_n 0.00421738f $X=7.51 $Y=2.465 $X2=0
+ $Y2=0
cc_545 N_A_398_74#_c_359_n N_VPWR_c_1657_n 0.0511446f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_546 N_A_398_74#_c_360_n N_VPWR_c_1657_n 0.00971754f $X=2.355 $Y=2.99 $X2=0
+ $Y2=0
cc_547 N_A_398_74#_c_367_n N_VPWR_c_1657_n 0.025655f $X=5.37 $Y=2.99 $X2=0 $Y2=0
cc_548 N_A_398_74#_c_368_n N_VPWR_c_1657_n 0.00583135f $X=4.78 $Y=2.99 $X2=0
+ $Y2=0
cc_549 N_A_398_74#_c_364_n A_728_463# 0.00497225f $X=3.79 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_550 N_A_398_74#_c_372_n A_1254_341# 0.00852216f $X=6.435 $Y=1.705 $X2=-0.19
+ $Y2=-0.245
cc_551 N_A_398_74#_c_340_n N_VGND_c_1856_n 0.0110038f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_552 N_A_398_74#_M1022_g N_VGND_c_1857_n 0.00147934f $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_553 N_A_398_74#_c_344_n N_VGND_c_1858_n 0.0287935f $X=6.52 $Y=1.12 $X2=0
+ $Y2=0
cc_554 N_A_398_74#_c_347_n N_VGND_c_1858_n 0.0106465f $X=6.605 $Y=0.34 $X2=0
+ $Y2=0
cc_555 N_A_398_74#_c_353_n N_VGND_c_1858_n 4.05806e-19 $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_556 N_A_398_74#_M1022_g N_VGND_c_1861_n 0.00527282f $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_557 N_A_398_74#_c_339_n N_VGND_c_1861_n 0.0591538f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_558 N_A_398_74#_c_340_n N_VGND_c_1861_n 0.0179217f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_559 N_A_398_74#_c_346_n N_VGND_c_1867_n 0.0617884f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_560 N_A_398_74#_c_347_n N_VGND_c_1867_n 0.0121867f $X=6.605 $Y=0.34 $X2=0
+ $Y2=0
cc_561 N_A_398_74#_c_353_n N_VGND_c_1867_n 0.00278271f $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_562 N_A_398_74#_M1022_g N_VGND_c_1870_n 0.00534666f $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_563 N_A_398_74#_c_339_n N_VGND_c_1870_n 0.0340476f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_564 N_A_398_74#_c_340_n N_VGND_c_1870_n 0.00971942f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_565 N_A_398_74#_c_346_n N_VGND_c_1870_n 0.0347045f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_566 N_A_398_74#_c_347_n N_VGND_c_1870_n 0.00660921f $X=6.605 $Y=0.34 $X2=0
+ $Y2=0
cc_567 N_A_398_74#_c_353_n N_VGND_c_1870_n 0.0035485f $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_568 N_A_398_74#_c_346_n N_VGND_c_1874_n 0.00587652f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_569 N_A_398_74#_c_351_n N_VGND_c_1874_n 0.00763101f $X=7.395 $Y=2.02 $X2=0
+ $Y2=0
cc_570 N_A_398_74#_c_344_n A_1262_74# 0.00897986f $X=6.52 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_571 N_A_398_74#_c_347_n A_1262_74# 6.58104e-19 $X=6.605 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_572 N_A_398_74#_c_346_n A_1462_74# 8.39422e-19 $X=7.39 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_573 N_A_398_74#_c_351_n A_1462_74# 0.0034631f $X=7.395 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_574 N_A_779_380#_c_641_n N_A_596_81#_c_740_n 0.017338f $X=4.95 $Y=1.885 $X2=0
+ $Y2=0
cc_575 N_A_779_380#_c_642_n N_A_596_81#_c_740_n 0.0139263f $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_576 N_A_779_380#_c_643_n N_A_596_81#_c_740_n 0.00677269f $X=5.115 $Y=2.515
+ $X2=0 $Y2=0
cc_577 N_A_779_380#_c_643_n N_A_596_81#_c_741_n 0.00895271f $X=5.115 $Y=2.515
+ $X2=0 $Y2=0
cc_578 N_A_779_380#_c_635_n N_A_596_81#_M1018_g 0.0153755f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_579 N_A_779_380#_c_637_n N_A_596_81#_M1018_g 0.00296272f $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_580 N_A_779_380#_c_641_n N_A_596_81#_c_727_n 0.0036927f $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_581 N_A_779_380#_c_635_n N_A_596_81#_c_727_n 7.42277e-19 $X=5.015 $Y=0.6
+ $X2=0 $Y2=0
cc_582 N_A_779_380#_c_636_n N_A_596_81#_c_727_n 0.0139263f $X=4.395 $Y=1.72
+ $X2=0 $Y2=0
cc_583 N_A_779_380#_c_632_n N_A_596_81#_c_728_n 0.00177919f $X=4.055 $Y=0.935
+ $X2=0 $Y2=0
cc_584 N_A_779_380#_c_632_n N_A_596_81#_c_729_n 0.0077045f $X=4.055 $Y=0.935
+ $X2=0 $Y2=0
cc_585 N_A_779_380#_c_633_n N_A_596_81#_c_729_n 0.00578861f $X=4.41 $Y=1.01
+ $X2=0 $Y2=0
cc_586 N_A_779_380#_c_634_n N_A_596_81#_c_729_n 0.00761441f $X=4.13 $Y=1.01
+ $X2=0 $Y2=0
cc_587 N_A_779_380#_c_635_n N_A_596_81#_c_729_n 0.0140413f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_588 N_A_779_380#_c_633_n N_A_596_81#_c_730_n 0.00406612f $X=4.41 $Y=1.01
+ $X2=0 $Y2=0
cc_589 N_A_779_380#_c_634_n N_A_596_81#_c_730_n 8.23249e-19 $X=4.13 $Y=1.01
+ $X2=0 $Y2=0
cc_590 N_A_779_380#_c_635_n N_A_596_81#_c_730_n 0.0156766f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_591 N_A_779_380#_c_637_n N_A_596_81#_c_730_n 0.00444456f $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_592 N_A_779_380#_c_633_n N_A_596_81#_c_731_n 0.00237419f $X=4.41 $Y=1.01
+ $X2=0 $Y2=0
cc_593 N_A_779_380#_c_641_n N_A_596_81#_c_731_n 0.0704401f $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_594 N_A_779_380#_c_642_n N_A_596_81#_c_731_n 0.00140465f $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_595 N_A_779_380#_c_635_n N_A_596_81#_c_731_n 0.0310993f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_596 N_A_779_380#_c_636_n N_A_596_81#_c_731_n 0.0123136f $X=4.395 $Y=1.72
+ $X2=0 $Y2=0
cc_597 N_A_779_380#_c_637_n N_A_596_81#_c_731_n 0.00126891f $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_598 N_A_779_380#_c_639_n N_A_596_81#_c_732_n 0.00247902f $X=4.23 $Y=1.975
+ $X2=0 $Y2=0
cc_599 N_A_779_380#_c_641_n N_A_596_81#_c_732_n 0.00453512f $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_600 N_A_779_380#_c_642_n N_A_596_81#_c_732_n 6.72497e-19 $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_601 N_A_779_380#_c_635_n N_A_596_81#_c_733_n 0.0363901f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_602 N_A_779_380#_c_637_n N_A_596_81#_c_733_n 2.43226e-19 $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_603 N_A_779_380#_c_636_n N_A_596_81#_c_734_n 5.72749e-19 $X=4.395 $Y=1.72
+ $X2=0 $Y2=0
cc_604 N_A_779_380#_c_640_n N_A_596_81#_c_736_n 9.56258e-19 $X=3.985 $Y=1.975
+ $X2=0 $Y2=0
cc_605 N_A_779_380#_c_641_n N_A_596_81#_c_739_n 4.77624e-19 $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_606 N_A_779_380#_c_635_n N_A_596_81#_c_739_n 0.00223707f $X=5.015 $Y=0.6
+ $X2=0 $Y2=0
cc_607 N_A_779_380#_c_636_n N_A_596_81#_c_739_n 0.00869085f $X=4.395 $Y=1.72
+ $X2=0 $Y2=0
cc_608 N_A_779_380#_c_637_n N_A_596_81#_c_739_n 0.0136391f $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_609 N_A_779_380#_c_643_n N_SET_B_c_896_n 0.00252974f $X=5.115 $Y=2.515 $X2=0
+ $Y2=0
cc_610 N_A_779_380#_c_643_n N_SET_B_c_897_n 0.00354543f $X=5.115 $Y=2.515 $X2=0
+ $Y2=0
cc_611 N_A_779_380#_c_635_n N_SET_B_M1028_g 0.00137951f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_612 N_A_779_380#_c_641_n N_SET_B_c_892_n 0.0129984f $X=4.95 $Y=1.885 $X2=0
+ $Y2=0
cc_613 N_A_779_380#_c_641_n N_SET_B_c_905_n 0.00232552f $X=4.95 $Y=1.885 $X2=0
+ $Y2=0
cc_614 N_A_779_380#_c_638_n N_A_225_74#_c_1049_n 0.00222169f $X=3.985 $Y=2.24
+ $X2=0 $Y2=0
cc_615 N_A_779_380#_c_638_n N_A_225_74#_c_1051_n 0.0214261f $X=3.985 $Y=2.24
+ $X2=0 $Y2=0
cc_616 N_A_779_380#_c_640_n N_A_225_74#_c_1051_n 0.00249329f $X=3.985 $Y=1.975
+ $X2=0 $Y2=0
cc_617 N_A_779_380#_c_638_n N_A_225_74#_c_1052_n 0.0103562f $X=3.985 $Y=2.24
+ $X2=0 $Y2=0
cc_618 N_A_779_380#_c_638_n N_VPWR_c_1660_n 0.00645065f $X=3.985 $Y=2.24 $X2=0
+ $Y2=0
cc_619 N_A_779_380#_c_638_n N_VPWR_c_1657_n 8.51577e-19 $X=3.985 $Y=2.24 $X2=0
+ $Y2=0
cc_620 N_A_779_380#_c_632_n N_VGND_c_1857_n 0.0108567f $X=4.055 $Y=0.935 $X2=0
+ $Y2=0
cc_621 N_A_779_380#_c_633_n N_VGND_c_1857_n 0.00687895f $X=4.41 $Y=1.01 $X2=0
+ $Y2=0
cc_622 N_A_779_380#_c_635_n N_VGND_c_1857_n 0.0244437f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_623 N_A_779_380#_c_635_n N_VGND_c_1858_n 0.0122754f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_624 N_A_779_380#_c_632_n N_VGND_c_1861_n 0.0045897f $X=4.055 $Y=0.935 $X2=0
+ $Y2=0
cc_625 N_A_779_380#_c_635_n N_VGND_c_1866_n 0.0175574f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_626 N_A_779_380#_c_632_n N_VGND_c_1870_n 0.0044912f $X=4.055 $Y=0.935 $X2=0
+ $Y2=0
cc_627 N_A_779_380#_c_635_n N_VGND_c_1870_n 0.019759f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_628 N_A_596_81#_c_741_n N_SET_B_c_896_n 0.00884898f $X=4.89 $Y=2.24 $X2=0
+ $Y2=0
cc_629 N_A_596_81#_c_725_n N_SET_B_c_896_n 0.0031279f $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_630 N_A_596_81#_c_741_n N_SET_B_c_897_n 0.0116352f $X=4.89 $Y=2.24 $X2=0
+ $Y2=0
cc_631 N_A_596_81#_c_725_n N_SET_B_c_897_n 0.00658537f $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_632 N_A_596_81#_c_723_n N_SET_B_M1028_g 0.00527452f $X=5.025 $Y=1.57 $X2=0
+ $Y2=0
cc_633 N_A_596_81#_M1018_g N_SET_B_M1028_g 0.0611842f $X=5.23 $Y=0.58 $X2=0
+ $Y2=0
cc_634 N_A_596_81#_c_725_n N_SET_B_M1028_g 0.0244411f $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_635 N_A_596_81#_c_726_n N_SET_B_M1028_g 0.0118733f $X=6.235 $Y=1.12 $X2=0
+ $Y2=0
cc_636 N_A_596_81#_c_731_n N_SET_B_M1028_g 0.00301751f $X=4.95 $Y=1.52 $X2=0
+ $Y2=0
cc_637 N_A_596_81#_c_733_n N_SET_B_M1028_g 3.61773e-19 $X=5.092 $Y=1.29 $X2=0
+ $Y2=0
cc_638 N_A_596_81#_c_734_n N_SET_B_M1028_g 0.00154129f $X=5.092 $Y=1.435 $X2=0
+ $Y2=0
cc_639 N_A_596_81#_c_735_n N_SET_B_M1028_g 0.0148959f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_640 N_A_596_81#_c_738_n N_SET_B_M1028_g 0.00115306f $X=6.1 $Y=1.205 $X2=0
+ $Y2=0
cc_641 N_A_596_81#_c_725_n N_SET_B_c_890_n 0.00355989f $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_642 N_A_596_81#_c_735_n N_SET_B_c_890_n 0.00860328f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_643 N_A_596_81#_c_738_n N_SET_B_c_890_n 0.00789782f $X=6.1 $Y=1.205 $X2=0
+ $Y2=0
cc_644 N_A_596_81#_c_740_n N_SET_B_c_891_n 2.72666e-19 $X=4.89 $Y=2.15 $X2=0
+ $Y2=0
cc_645 N_A_596_81#_c_727_n N_SET_B_c_891_n 9.05772e-19 $X=5.025 $Y=1.645 $X2=0
+ $Y2=0
cc_646 N_A_596_81#_c_731_n N_SET_B_c_891_n 0.00172913f $X=4.95 $Y=1.52 $X2=0
+ $Y2=0
cc_647 N_A_596_81#_c_735_n N_SET_B_c_891_n 0.00314092f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_648 N_A_596_81#_c_740_n N_SET_B_c_892_n 6.13227e-19 $X=4.89 $Y=2.15 $X2=0
+ $Y2=0
cc_649 N_A_596_81#_c_725_n N_SET_B_c_892_n 7.06984e-19 $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_650 N_A_596_81#_c_727_n N_SET_B_c_892_n 0.00124776f $X=5.025 $Y=1.645 $X2=0
+ $Y2=0
cc_651 N_A_596_81#_c_731_n N_SET_B_c_892_n 0.00404118f $X=4.95 $Y=1.52 $X2=0
+ $Y2=0
cc_652 N_A_596_81#_c_735_n N_SET_B_c_892_n 0.0119231f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_653 N_A_596_81#_c_740_n N_SET_B_c_905_n 0.00884898f $X=4.89 $Y=2.15 $X2=0
+ $Y2=0
cc_654 N_A_596_81#_c_725_n N_SET_B_c_905_n 0.00769918f $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_655 N_A_596_81#_c_727_n N_SET_B_c_905_n 0.0065664f $X=5.025 $Y=1.645 $X2=0
+ $Y2=0
cc_656 N_A_596_81#_c_735_n N_SET_B_c_905_n 0.00384007f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_657 N_A_596_81#_c_728_n N_A_225_74#_M1008_g 8.37131e-19 $X=3.45 $Y=0.615
+ $X2=0 $Y2=0
cc_658 N_A_596_81#_c_744_n N_A_225_74#_c_1051_n 0.00627699f $X=3.34 $Y=2.515
+ $X2=0 $Y2=0
cc_659 N_A_596_81#_c_736_n N_A_225_74#_c_1051_n 0.00292835f $X=3.355 $Y=2.295
+ $X2=0 $Y2=0
cc_660 N_A_596_81#_c_741_n N_A_225_74#_c_1052_n 0.00882199f $X=4.89 $Y=2.24
+ $X2=0 $Y2=0
cc_661 N_A_596_81#_c_725_n N_A_225_74#_c_1052_n 0.00907339f $X=6.195 $Y=1.63
+ $X2=0 $Y2=0
cc_662 N_A_596_81#_c_725_n N_A_225_74#_M1013_g 0.0330539f $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_663 N_A_596_81#_c_725_n N_A_225_74#_c_1038_n 0.00553621f $X=6.195 $Y=1.63
+ $X2=0 $Y2=0
cc_664 N_A_596_81#_c_725_n N_A_1355_377#_c_1366_n 0.00183199f $X=6.195 $Y=1.63
+ $X2=0 $Y2=0
cc_665 N_A_596_81#_c_725_n N_A_1355_377#_c_1355_n 0.0016321f $X=6.195 $Y=1.63
+ $X2=0 $Y2=0
cc_666 N_A_596_81#_c_725_n N_A_1355_377#_c_1360_n 7.49332e-19 $X=6.195 $Y=1.63
+ $X2=0 $Y2=0
cc_667 N_A_596_81#_c_744_n N_A_27_80#_c_1597_n 0.0183821f $X=3.34 $Y=2.515 $X2=0
+ $Y2=0
cc_668 N_A_596_81#_c_736_n N_A_27_80#_c_1597_n 0.00583359f $X=3.355 $Y=2.295
+ $X2=0 $Y2=0
cc_669 N_A_596_81#_c_725_n N_VPWR_c_1661_n 0.0113891f $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_670 N_A_596_81#_c_725_n N_VPWR_c_1657_n 9.49986e-19 $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_671 N_A_596_81#_c_728_n N_VGND_c_1857_n 0.0102369f $X=3.45 $Y=0.615 $X2=0
+ $Y2=0
cc_672 N_A_596_81#_c_729_n N_VGND_c_1857_n 0.0136266f $X=4.115 $Y=0.97 $X2=0
+ $Y2=0
cc_673 N_A_596_81#_c_725_n N_VGND_c_1858_n 0.00159559f $X=6.195 $Y=1.63 $X2=0
+ $Y2=0
cc_674 N_A_596_81#_c_726_n N_VGND_c_1858_n 0.0113166f $X=6.235 $Y=1.12 $X2=0
+ $Y2=0
cc_675 N_A_596_81#_c_735_n N_VGND_c_1858_n 0.00656613f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_676 N_A_596_81#_c_738_n N_VGND_c_1858_n 0.0179048f $X=6.1 $Y=1.205 $X2=0
+ $Y2=0
cc_677 N_A_596_81#_c_728_n N_VGND_c_1861_n 0.00962837f $X=3.45 $Y=0.615 $X2=0
+ $Y2=0
cc_678 N_A_596_81#_M1018_g N_VGND_c_1866_n 0.00434997f $X=5.23 $Y=0.58 $X2=0
+ $Y2=0
cc_679 N_A_596_81#_c_726_n N_VGND_c_1867_n 0.00383152f $X=6.235 $Y=1.12 $X2=0
+ $Y2=0
cc_680 N_A_596_81#_M1018_g N_VGND_c_1870_n 0.00824278f $X=5.23 $Y=0.58 $X2=0
+ $Y2=0
cc_681 N_A_596_81#_c_726_n N_VGND_c_1870_n 0.00758168f $X=6.235 $Y=1.12 $X2=0
+ $Y2=0
cc_682 N_A_596_81#_c_728_n N_VGND_c_1870_n 0.00894094f $X=3.45 $Y=0.615 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_897_n N_A_225_74#_c_1052_n 0.00946336f $X=5.4 $Y=2.24 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_890_n N_A_225_74#_c_1037_n 0.00355894f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_890_n N_A_225_74#_c_1038_n 0.00690366f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_890_n N_A_225_74#_M1032_g 0.00409351f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_687 N_SET_B_M1025_g N_A_1510_48#_M1030_g 0.0563813f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_894_n N_A_1510_48#_M1030_g 0.00223551f $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_889_n N_A_1510_48#_c_1222_n 0.0247275f $X=8.415 $Y=2.155 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_899_n N_A_1510_48#_c_1223_n 0.00998154f $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_691 N_SET_B_M1025_g N_A_1510_48#_c_1214_n 0.00739584f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_887_n N_A_1510_48#_c_1214_n 0.00256307f $X=8.34 $Y=1.3 $X2=0
+ $Y2=0
cc_693 N_SET_B_c_888_n N_A_1510_48#_c_1214_n 0.00453006f $X=8.09 $Y=1.3 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_889_n N_A_1510_48#_c_1214_n 9.56134e-19 $X=8.415 $Y=2.155 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_890_n N_A_1510_48#_c_1214_n 0.025713f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_696 SET_B N_A_1510_48#_c_1214_n 0.00265164f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_697 N_SET_B_c_894_n N_A_1510_48#_c_1214_n 8.16272e-19 $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_698 N_SET_B_c_895_n N_A_1510_48#_c_1214_n 0.0424843f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_699 N_SET_B_c_887_n N_A_1510_48#_c_1215_n 0.0084215f $X=8.34 $Y=1.3 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_890_n N_A_1510_48#_c_1215_n 0.00472787f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_701 SET_B N_A_1510_48#_c_1215_n 0.00196951f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_702 N_SET_B_c_895_n N_A_1510_48#_c_1215_n 0.031422f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_703 N_SET_B_M1025_g N_A_1510_48#_c_1216_n 0.0108479f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_704 N_SET_B_c_899_n N_A_1510_48#_c_1224_n 7.90532e-19 $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_899_n N_A_1510_48#_c_1226_n 3.94558e-19 $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_889_n N_A_1510_48#_c_1226_n 3.21135e-19 $X=8.415 $Y=2.155 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_888_n N_A_1510_48#_c_1221_n 0.0104108f $X=8.09 $Y=1.3 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_889_n N_A_1510_48#_c_1221_n 0.0188382f $X=8.415 $Y=2.155 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_890_n N_A_1510_48#_c_1221_n 0.0105411f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_710 SET_B N_A_1510_48#_c_1221_n 8.64502e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_711 N_SET_B_c_895_n N_A_1510_48#_c_1221_n 9.42269e-19 $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_712 N_SET_B_M1025_g N_A_1355_377#_c_1334_n 0.00678433f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_895_n N_A_1355_377#_c_1335_n 0.00122225f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_889_n N_A_1355_377#_c_1339_n 0.0124328f $X=8.415 $Y=2.155 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_894_n N_A_1355_377#_c_1339_n 0.0101337f $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_895_n N_A_1355_377#_c_1339_n 0.00368499f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_717 N_SET_B_c_890_n N_A_1355_377#_c_1344_n 0.0130228f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_718 N_SET_B_c_887_n N_A_1355_377#_c_1356_n 0.00442681f $X=8.34 $Y=1.3 $X2=0
+ $Y2=0
cc_719 N_SET_B_c_899_n N_A_1355_377#_c_1356_n 0.00378805f $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_720 N_SET_B_c_889_n N_A_1355_377#_c_1356_n 0.0129397f $X=8.415 $Y=2.155 $X2=0
+ $Y2=0
cc_721 N_SET_B_c_890_n N_A_1355_377#_c_1356_n 0.00672574f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_722 SET_B N_A_1355_377#_c_1356_n 0.00261165f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_723 N_SET_B_c_895_n N_A_1355_377#_c_1356_n 0.00628568f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_899_n N_A_1355_377#_c_1357_n 0.00857431f $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_889_n N_A_1355_377#_c_1345_n 0.00158354f $X=8.415 $Y=2.155
+ $X2=0 $Y2=0
cc_726 SET_B N_A_1355_377#_c_1345_n 0.00118411f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_727 N_SET_B_c_894_n N_A_1355_377#_c_1345_n 0.00149353f $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_728 N_SET_B_c_895_n N_A_1355_377#_c_1345_n 0.0216237f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_729 N_SET_B_c_890_n N_A_1355_377#_c_1360_n 0.0266747f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_730 N_SET_B_c_899_n N_A_1355_377#_c_1363_n 4.54623e-19 $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_731 N_SET_B_c_890_n N_A_1355_377#_c_1363_n 0.00355761f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_732 N_SET_B_c_899_n N_A_1355_377#_c_1364_n 2.84963e-19 $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_889_n N_A_1355_377#_c_1364_n 0.0114654f $X=8.415 $Y=2.155 $X2=0
+ $Y2=0
cc_734 SET_B N_A_1355_377#_c_1364_n 8.38169e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_735 N_SET_B_c_894_n N_A_1355_377#_c_1364_n 8.70886e-19 $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_736 N_SET_B_c_895_n N_A_1355_377#_c_1364_n 0.0129183f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_737 N_SET_B_c_897_n N_VPWR_c_1661_n 0.00160015f $X=5.4 $Y=2.24 $X2=0 $Y2=0
cc_738 N_SET_B_c_899_n N_VPWR_c_1662_n 0.00373065f $X=8.38 $Y=2.465 $X2=0 $Y2=0
cc_739 N_SET_B_c_899_n N_VPWR_c_1671_n 0.00445602f $X=8.38 $Y=2.465 $X2=0 $Y2=0
cc_740 N_SET_B_c_899_n N_VPWR_c_1657_n 0.00459843f $X=8.38 $Y=2.465 $X2=0 $Y2=0
cc_741 N_SET_B_M1028_g N_VGND_c_1858_n 0.0128389f $X=5.62 $Y=0.58 $X2=0 $Y2=0
cc_742 N_SET_B_M1028_g N_VGND_c_1866_n 0.00461464f $X=5.62 $Y=0.58 $X2=0 $Y2=0
cc_743 N_SET_B_M1025_g N_VGND_c_1867_n 0.00384553f $X=8.015 $Y=0.58 $X2=0 $Y2=0
cc_744 N_SET_B_M1028_g N_VGND_c_1870_n 0.00910593f $X=5.62 $Y=0.58 $X2=0 $Y2=0
cc_745 N_SET_B_M1025_g N_VGND_c_1870_n 0.00383468f $X=8.015 $Y=0.58 $X2=0 $Y2=0
cc_746 N_SET_B_M1025_g N_VGND_c_1874_n 0.0107673f $X=8.015 $Y=0.58 $X2=0 $Y2=0
cc_747 N_SET_B_c_887_n N_VGND_c_1874_n 2.20993e-19 $X=8.34 $Y=1.3 $X2=0 $Y2=0
cc_748 N_A_225_74#_M1032_g N_A_1510_48#_M1030_g 0.0378389f $X=7.235 $Y=0.58
+ $X2=0 $Y2=0
cc_749 N_A_225_74#_c_1037_n N_A_1510_48#_c_1221_n 0.039364f $X=7.16 $Y=1.735
+ $X2=0 $Y2=0
cc_750 N_A_225_74#_M1013_g N_A_1355_377#_c_1366_n 0.00747649f $X=6.7 $Y=2.385
+ $X2=0 $Y2=0
cc_751 N_A_225_74#_c_1037_n N_A_1355_377#_c_1354_n 0.00139562f $X=7.16 $Y=1.735
+ $X2=0 $Y2=0
cc_752 N_A_225_74#_M1013_g N_A_1355_377#_c_1355_n 0.012333f $X=6.7 $Y=2.385
+ $X2=0 $Y2=0
cc_753 N_A_225_74#_c_1059_n N_A_1355_377#_c_1355_n 4.34896e-19 $X=6.7 $Y=3.15
+ $X2=0 $Y2=0
cc_754 N_A_225_74#_c_1037_n N_A_1355_377#_c_1344_n 0.00327799f $X=7.16 $Y=1.735
+ $X2=0 $Y2=0
cc_755 N_A_225_74#_M1032_g N_A_1355_377#_c_1344_n 0.0162403f $X=7.235 $Y=0.58
+ $X2=0 $Y2=0
cc_756 N_A_225_74#_M1013_g N_A_1355_377#_c_1360_n 0.0101622f $X=6.7 $Y=2.385
+ $X2=0 $Y2=0
cc_757 N_A_225_74#_c_1037_n N_A_1355_377#_c_1360_n 0.0182349f $X=7.16 $Y=1.735
+ $X2=0 $Y2=0
cc_758 N_A_225_74#_M1032_g N_A_1355_377#_c_1346_n 0.00979462f $X=7.235 $Y=0.58
+ $X2=0 $Y2=0
cc_759 N_A_225_74#_M1027_s N_A_27_80#_c_1596_n 0.0126187f $X=1.145 $Y=1.79 $X2=0
+ $Y2=0
cc_760 N_A_225_74#_c_1061_n N_A_27_80#_c_1596_n 0.0190006f $X=1.305 $Y=1.87
+ $X2=0 $Y2=0
cc_761 N_A_225_74#_c_1062_n N_A_27_80#_c_1596_n 0.0142272f $X=1.145 $Y=1.87
+ $X2=0 $Y2=0
cc_762 N_A_225_74#_c_1063_n N_A_27_80#_c_1596_n 0.0057885f $X=2.025 $Y=1.805
+ $X2=0 $Y2=0
cc_763 N_A_225_74#_c_1034_n N_A_27_80#_c_1597_n 0.0150147f $X=1.965 $Y=1.715
+ $X2=0 $Y2=0
cc_764 N_A_225_74#_c_1046_n N_A_27_80#_c_1597_n 0.0301029f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_765 N_A_225_74#_c_1041_n N_A_27_80#_c_1597_n 0.00284892f $X=2.41 $Y=1.465
+ $X2=0 $Y2=0
cc_766 N_A_225_74#_c_1063_n N_A_27_80#_c_1597_n 0.0337756f $X=2.025 $Y=1.805
+ $X2=0 $Y2=0
cc_767 N_A_225_74#_M1017_g N_A_27_80#_c_1591_n 8.15758e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_768 N_A_225_74#_c_1034_n N_A_27_80#_c_1591_n 0.00100001f $X=1.965 $Y=1.715
+ $X2=0 $Y2=0
cc_769 N_A_225_74#_c_1046_n N_A_27_80#_c_1591_n 0.00931709f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_770 N_A_225_74#_c_1035_n N_A_27_80#_c_1591_n 0.0104106f $X=2.83 $Y=1.12 $X2=0
+ $Y2=0
cc_771 N_A_225_74#_M1008_g N_A_27_80#_c_1591_n 0.00434152f $X=2.905 $Y=0.615
+ $X2=0 $Y2=0
cc_772 N_A_225_74#_c_1040_n N_A_27_80#_c_1591_n 0.0147929f $X=2.485 $Y=1.12
+ $X2=0 $Y2=0
cc_773 N_A_225_74#_c_1063_n N_A_27_80#_c_1591_n 0.0137141f $X=2.025 $Y=1.805
+ $X2=0 $Y2=0
cc_774 N_A_225_74#_c_1043_n N_A_27_80#_c_1591_n 0.0302853f $X=2.19 $Y=1.465
+ $X2=0 $Y2=0
cc_775 N_A_225_74#_c_1034_n N_A_27_80#_c_1641_n 0.00326455f $X=1.965 $Y=1.715
+ $X2=0 $Y2=0
cc_776 N_A_225_74#_c_1063_n N_A_27_80#_c_1641_n 0.0112057f $X=2.025 $Y=1.805
+ $X2=0 $Y2=0
cc_777 N_A_225_74#_c_1035_n N_A_27_80#_c_1593_n 0.00467868f $X=2.83 $Y=1.12
+ $X2=0 $Y2=0
cc_778 N_A_225_74#_M1008_g N_A_27_80#_c_1593_n 0.00437989f $X=2.905 $Y=0.615
+ $X2=0 $Y2=0
cc_779 N_A_225_74#_c_1063_n N_VPWR_M1027_d 0.00196757f $X=2.025 $Y=1.805 $X2=0
+ $Y2=0
cc_780 N_A_225_74#_c_1034_n N_VPWR_c_1659_n 0.00764723f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_781 N_A_225_74#_c_1046_n N_VPWR_c_1659_n 3.21585e-19 $X=2.485 $Y=3.075 $X2=0
+ $Y2=0
cc_782 N_A_225_74#_c_1048_n N_VPWR_c_1659_n 0.00272925f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_783 N_A_225_74#_c_1050_n N_VPWR_c_1660_n 8.5651e-19 $X=3.565 $Y=3.075 $X2=0
+ $Y2=0
cc_784 N_A_225_74#_c_1052_n N_VPWR_c_1660_n 0.0292393f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_785 N_A_225_74#_c_1052_n N_VPWR_c_1661_n 0.0264687f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_786 N_A_225_74#_M1013_g N_VPWR_c_1661_n 0.00378611f $X=6.7 $Y=2.385 $X2=0
+ $Y2=0
cc_787 N_A_225_74#_c_1059_n N_VPWR_c_1661_n 0.00290668f $X=6.7 $Y=3.15 $X2=0
+ $Y2=0
cc_788 N_A_225_74#_c_1052_n N_VPWR_c_1665_n 0.0262935f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_789 N_A_225_74#_c_1034_n N_VPWR_c_1669_n 0.0048608f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_790 N_A_225_74#_c_1048_n N_VPWR_c_1669_n 0.0372724f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_791 N_A_225_74#_c_1052_n N_VPWR_c_1670_n 0.0306837f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_792 N_A_225_74#_c_1034_n N_VPWR_c_1657_n 0.00480464f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_793 N_A_225_74#_c_1047_n N_VPWR_c_1657_n 0.0215278f $X=3.475 $Y=3.15 $X2=0
+ $Y2=0
cc_794 N_A_225_74#_c_1048_n N_VPWR_c_1657_n 0.00604517f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_795 N_A_225_74#_c_1052_n N_VPWR_c_1657_n 0.0779542f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_796 N_A_225_74#_c_1058_n N_VPWR_c_1657_n 0.00441524f $X=3.565 $Y=3.15 $X2=0
+ $Y2=0
cc_797 N_A_225_74#_c_1059_n N_VPWR_c_1657_n 0.0122301f $X=6.7 $Y=3.15 $X2=0
+ $Y2=0
cc_798 N_A_225_74#_c_1044_n N_VGND_c_1854_n 0.0387749f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_799 N_A_225_74#_c_1044_n N_VGND_c_1855_n 0.0203368f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_800 N_A_225_74#_M1017_g N_VGND_c_1856_n 0.0115714f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_801 N_A_225_74#_c_1044_n N_VGND_c_1856_n 0.0268179f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_802 N_A_225_74#_M1017_g N_VGND_c_1861_n 0.00383152f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_803 N_A_225_74#_M1008_g N_VGND_c_1861_n 9.15902e-19 $X=2.905 $Y=0.615 $X2=0
+ $Y2=0
cc_804 N_A_225_74#_M1032_g N_VGND_c_1867_n 0.00278271f $X=7.235 $Y=0.58 $X2=0
+ $Y2=0
cc_805 N_A_225_74#_M1017_g N_VGND_c_1870_n 0.00762539f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_806 N_A_225_74#_M1032_g N_VGND_c_1870_n 0.00353931f $X=7.235 $Y=0.58 $X2=0
+ $Y2=0
cc_807 N_A_225_74#_c_1044_n N_VGND_c_1870_n 0.0167889f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_808 N_A_1510_48#_c_1215_n N_A_1355_377#_c_1334_n 0.00361072f $X=8.925
+ $Y=0.925 $X2=0 $Y2=0
cc_809 N_A_1510_48#_c_1217_n N_A_1355_377#_c_1334_n 0.0116357f $X=9.09 $Y=0.58
+ $X2=0 $Y2=0
cc_810 N_A_1510_48#_c_1220_n N_A_1355_377#_c_1334_n 6.34661e-19 $X=9.09 $Y=0.925
+ $X2=0 $Y2=0
cc_811 N_A_1510_48#_c_1219_n N_A_1355_377#_c_1336_n 0.00619224f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_812 N_A_1510_48#_c_1224_n N_A_1355_377#_c_1348_n 0.0127509f $X=9.165 $Y=2.75
+ $X2=0 $Y2=0
cc_813 N_A_1510_48#_c_1225_n N_A_1355_377#_c_1348_n 0.0192416f $X=9.565 $Y=2.475
+ $X2=0 $Y2=0
cc_814 N_A_1510_48#_c_1226_n N_A_1355_377#_c_1348_n 0.00203684f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_815 N_A_1510_48#_c_1219_n N_A_1355_377#_c_1348_n 0.00451981f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_816 N_A_1510_48#_c_1217_n N_A_1355_377#_c_1337_n 0.0043971f $X=9.09 $Y=0.58
+ $X2=0 $Y2=0
cc_817 N_A_1510_48#_c_1218_n N_A_1355_377#_c_1337_n 0.00231095f $X=9.565
+ $Y=0.925 $X2=0 $Y2=0
cc_818 N_A_1510_48#_c_1219_n N_A_1355_377#_c_1337_n 0.00225427f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_819 N_A_1510_48#_c_1225_n N_A_1355_377#_c_1349_n 0.00176747f $X=9.565
+ $Y=2.475 $X2=0 $Y2=0
cc_820 N_A_1510_48#_c_1219_n N_A_1355_377#_c_1349_n 0.0054501f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_821 N_A_1510_48#_c_1218_n N_A_1355_377#_c_1339_n 0.00736519f $X=9.565
+ $Y=0.925 $X2=0 $Y2=0
cc_822 N_A_1510_48#_c_1219_n N_A_1355_377#_c_1339_n 0.0294834f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_823 N_A_1510_48#_c_1215_n N_A_1355_377#_c_1342_n 0.00925086f $X=8.925
+ $Y=0.925 $X2=0 $Y2=0
cc_824 N_A_1510_48#_c_1219_n N_A_1355_377#_c_1342_n 0.00382379f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_825 N_A_1510_48#_c_1220_n N_A_1355_377#_c_1342_n 0.0207635f $X=9.09 $Y=0.925
+ $X2=0 $Y2=0
cc_826 N_A_1510_48#_M1030_g N_A_1355_377#_c_1344_n 6.67309e-19 $X=7.625 $Y=0.58
+ $X2=0 $Y2=0
cc_827 N_A_1510_48#_c_1222_n N_A_1355_377#_c_1356_n 0.00909196f $X=7.93 $Y=2.375
+ $X2=0 $Y2=0
cc_828 N_A_1510_48#_c_1223_n N_A_1355_377#_c_1356_n 0.00521664f $X=7.93 $Y=2.465
+ $X2=0 $Y2=0
cc_829 N_A_1510_48#_c_1221_n N_A_1355_377#_c_1356_n 0.0019319f $X=7.93 $Y=1.75
+ $X2=0 $Y2=0
cc_830 N_A_1510_48#_c_1223_n N_A_1355_377#_c_1357_n 5.32065e-19 $X=7.93 $Y=2.465
+ $X2=0 $Y2=0
cc_831 N_A_1510_48#_c_1224_n N_A_1355_377#_c_1357_n 0.0282824f $X=9.165 $Y=2.75
+ $X2=0 $Y2=0
cc_832 N_A_1510_48#_c_1226_n N_A_1355_377#_c_1357_n 0.00568938f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_833 N_A_1510_48#_c_1226_n N_A_1355_377#_c_1358_n 0.00538906f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_834 N_A_1510_48#_c_1225_n N_A_1355_377#_c_1359_n 0.00507721f $X=9.565
+ $Y=2.475 $X2=0 $Y2=0
cc_835 N_A_1510_48#_c_1226_n N_A_1355_377#_c_1359_n 0.0233648f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_836 N_A_1510_48#_c_1219_n N_A_1355_377#_c_1359_n 0.0135838f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_837 N_A_1510_48#_c_1218_n N_A_1355_377#_c_1345_n 0.00978752f $X=9.565
+ $Y=0.925 $X2=0 $Y2=0
cc_838 N_A_1510_48#_c_1219_n N_A_1355_377#_c_1345_n 0.0615164f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_839 N_A_1510_48#_c_1220_n N_A_1355_377#_c_1345_n 0.0140685f $X=9.09 $Y=0.925
+ $X2=0 $Y2=0
cc_840 N_A_1510_48#_M1030_g N_A_1355_377#_c_1346_n 2.73884e-19 $X=7.625 $Y=0.58
+ $X2=0 $Y2=0
cc_841 N_A_1510_48#_c_1223_n N_A_1355_377#_c_1361_n 7.54283e-19 $X=7.93 $Y=2.465
+ $X2=0 $Y2=0
cc_842 N_A_1510_48#_c_1222_n N_A_1355_377#_c_1363_n 0.00456539f $X=7.93 $Y=2.375
+ $X2=0 $Y2=0
cc_843 N_A_1510_48#_c_1223_n N_A_1355_377#_c_1363_n 0.00760762f $X=7.93 $Y=2.465
+ $X2=0 $Y2=0
cc_844 N_A_1510_48#_c_1214_n N_A_1355_377#_c_1363_n 0.0257755f $X=7.935 $Y=1.75
+ $X2=0 $Y2=0
cc_845 N_A_1510_48#_c_1221_n N_A_1355_377#_c_1363_n 0.00292111f $X=7.93 $Y=1.75
+ $X2=0 $Y2=0
cc_846 N_A_1510_48#_c_1226_n N_A_1355_377#_c_1364_n 0.00681171f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_847 N_A_1510_48#_c_1225_n N_VPWR_M1006_d 0.00346493f $X=9.565 $Y=2.475 $X2=0
+ $Y2=0
cc_848 N_A_1510_48#_c_1219_n N_VPWR_M1006_d 0.00837897f $X=9.65 $Y=2.39 $X2=0
+ $Y2=0
cc_849 N_A_1510_48#_c_1223_n N_VPWR_c_1662_n 0.00623994f $X=7.93 $Y=2.465 $X2=0
+ $Y2=0
cc_850 N_A_1510_48#_c_1224_n N_VPWR_c_1663_n 0.00869586f $X=9.165 $Y=2.75 $X2=0
+ $Y2=0
cc_851 N_A_1510_48#_c_1225_n N_VPWR_c_1663_n 0.0111424f $X=9.565 $Y=2.475 $X2=0
+ $Y2=0
cc_852 N_A_1510_48#_c_1223_n N_VPWR_c_1665_n 0.00422316f $X=7.93 $Y=2.465 $X2=0
+ $Y2=0
cc_853 N_A_1510_48#_c_1224_n N_VPWR_c_1671_n 0.0144853f $X=9.165 $Y=2.75 $X2=0
+ $Y2=0
cc_854 N_A_1510_48#_c_1223_n N_VPWR_c_1657_n 0.00453881f $X=7.93 $Y=2.465 $X2=0
+ $Y2=0
cc_855 N_A_1510_48#_c_1224_n N_VPWR_c_1657_n 0.0120561f $X=9.165 $Y=2.75 $X2=0
+ $Y2=0
cc_856 N_A_1510_48#_c_1225_n N_VPWR_c_1657_n 0.0080698f $X=9.565 $Y=2.475 $X2=0
+ $Y2=0
cc_857 N_A_1510_48#_c_1218_n N_Q_N_c_1803_n 0.00764487f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_858 N_A_1510_48#_c_1225_n Q_N 0.00787809f $X=9.565 $Y=2.475 $X2=0 $Y2=0
cc_859 N_A_1510_48#_c_1219_n Q_N 0.0432234f $X=9.65 $Y=2.39 $X2=0 $Y2=0
cc_860 N_A_1510_48#_c_1218_n N_Q_N_c_1805_n 0.00277175f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_861 N_A_1510_48#_c_1219_n N_Q_N_c_1805_n 0.0148084f $X=9.65 $Y=2.39 $X2=0
+ $Y2=0
cc_862 N_A_1510_48#_c_1218_n N_VGND_M1014_s 0.00702554f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_863 N_A_1510_48#_c_1219_n N_VGND_M1014_s 0.00245883f $X=9.65 $Y=2.39 $X2=0
+ $Y2=0
cc_864 N_A_1510_48#_c_1217_n N_VGND_c_1859_n 0.0171919f $X=9.09 $Y=0.58 $X2=0
+ $Y2=0
cc_865 N_A_1510_48#_c_1218_n N_VGND_c_1859_n 0.0212677f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_866 N_A_1510_48#_c_1217_n N_VGND_c_1863_n 0.0102067f $X=9.09 $Y=0.58 $X2=0
+ $Y2=0
cc_867 N_A_1510_48#_M1030_g N_VGND_c_1867_n 0.00449242f $X=7.625 $Y=0.58 $X2=0
+ $Y2=0
cc_868 N_A_1510_48#_M1030_g N_VGND_c_1870_n 0.00871678f $X=7.625 $Y=0.58 $X2=0
+ $Y2=0
cc_869 N_A_1510_48#_c_1215_n N_VGND_c_1870_n 0.00709649f $X=8.925 $Y=0.925 $X2=0
+ $Y2=0
cc_870 N_A_1510_48#_c_1216_n N_VGND_c_1870_n 0.0108158f $X=8.1 $Y=0.925 $X2=0
+ $Y2=0
cc_871 N_A_1510_48#_c_1217_n N_VGND_c_1870_n 0.0114381f $X=9.09 $Y=0.58 $X2=0
+ $Y2=0
cc_872 N_A_1510_48#_c_1218_n N_VGND_c_1870_n 0.00883761f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_873 N_A_1510_48#_M1030_g N_VGND_c_1874_n 0.00126877f $X=7.625 $Y=0.58 $X2=0
+ $Y2=0
cc_874 N_A_1510_48#_c_1215_n N_VGND_c_1874_n 0.0502316f $X=8.925 $Y=0.925 $X2=0
+ $Y2=0
cc_875 N_A_1510_48#_c_1216_n N_VGND_c_1874_n 0.00238625f $X=8.1 $Y=0.925 $X2=0
+ $Y2=0
cc_876 N_A_1355_377#_c_1341_n N_A_2113_74#_c_1534_n 7.26921e-19 $X=10.925
+ $Y=1.79 $X2=0 $Y2=0
cc_877 N_A_1355_377#_c_1352_n N_A_2113_74#_c_1534_n 0.0189706f $X=10.99 $Y=1.94
+ $X2=0 $Y2=0
cc_878 N_A_1355_377#_c_1343_n N_A_2113_74#_c_1534_n 0.0240488f $X=10.925 $Y=1.41
+ $X2=0 $Y2=0
cc_879 N_A_1355_377#_c_1353_n N_A_2113_74#_c_1534_n 0.00528982f $X=10.99
+ $Y=1.865 $X2=0 $Y2=0
cc_880 N_A_1355_377#_M1026_g N_A_2113_74#_c_1535_n 0.0205551f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_881 N_A_1355_377#_c_1337_n N_A_2113_74#_c_1536_n 0.00119747f $X=9.935 $Y=1.21
+ $X2=0 $Y2=0
cc_882 N_A_1355_377#_M1026_g N_A_2113_74#_c_1536_n 0.00674464f $X=10.925
+ $Y=0.645 $X2=0 $Y2=0
cc_883 N_A_1355_377#_c_1337_n N_A_2113_74#_c_1537_n 3.90625e-19 $X=9.935 $Y=1.21
+ $X2=0 $Y2=0
cc_884 N_A_1355_377#_c_1338_n N_A_2113_74#_c_1537_n 0.00224708f $X=10.85 $Y=1.41
+ $X2=0 $Y2=0
cc_885 N_A_1355_377#_M1026_g N_A_2113_74#_c_1537_n 0.0099886f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_886 N_A_1355_377#_c_1338_n N_A_2113_74#_c_1538_n 0.00711579f $X=10.85 $Y=1.41
+ $X2=0 $Y2=0
cc_887 N_A_1355_377#_c_1341_n N_A_2113_74#_c_1538_n 0.0138825f $X=10.925 $Y=1.79
+ $X2=0 $Y2=0
cc_888 N_A_1355_377#_c_1352_n N_A_2113_74#_c_1538_n 0.00865733f $X=10.99 $Y=1.94
+ $X2=0 $Y2=0
cc_889 N_A_1355_377#_c_1343_n N_A_2113_74#_c_1539_n 0.0191447f $X=10.925 $Y=1.41
+ $X2=0 $Y2=0
cc_890 N_A_1355_377#_c_1353_n N_A_2113_74#_c_1539_n 0.00279973f $X=10.99
+ $Y=1.865 $X2=0 $Y2=0
cc_891 N_A_1355_377#_c_1338_n N_A_2113_74#_c_1540_n 0.00533007f $X=10.85 $Y=1.41
+ $X2=0 $Y2=0
cc_892 N_A_1355_377#_M1026_g N_A_2113_74#_c_1540_n 0.00377159f $X=10.925
+ $Y=0.645 $X2=0 $Y2=0
cc_893 N_A_1355_377#_c_1338_n N_A_2113_74#_c_1560_n 0.0110675f $X=10.85 $Y=1.41
+ $X2=0 $Y2=0
cc_894 N_A_1355_377#_c_1343_n N_A_2113_74#_c_1560_n 0.00192549f $X=10.925
+ $Y=1.41 $X2=0 $Y2=0
cc_895 N_A_1355_377#_c_1356_n N_VPWR_c_1662_n 0.0145069f $X=8.44 $Y=2.265 $X2=0
+ $Y2=0
cc_896 N_A_1355_377#_c_1357_n N_VPWR_c_1662_n 0.0215225f $X=8.605 $Y=2.75 $X2=0
+ $Y2=0
cc_897 N_A_1355_377#_c_1361_n N_VPWR_c_1662_n 0.00712065f $X=7.45 $Y=2.692 $X2=0
+ $Y2=0
cc_898 N_A_1355_377#_c_1348_n N_VPWR_c_1663_n 0.00348428f $X=9.475 $Y=2.465
+ $X2=0 $Y2=0
cc_899 N_A_1355_377#_c_1349_n N_VPWR_c_1663_n 0.00873738f $X=9.98 $Y=1.765 $X2=0
+ $Y2=0
cc_900 N_A_1355_377#_c_1352_n N_VPWR_c_1664_n 0.0161758f $X=10.99 $Y=1.94 $X2=0
+ $Y2=0
cc_901 N_A_1355_377#_c_1353_n N_VPWR_c_1664_n 4.22058e-19 $X=10.99 $Y=1.865
+ $X2=0 $Y2=0
cc_902 N_A_1355_377#_c_1354_n N_VPWR_c_1665_n 0.0133586f $X=7.238 $Y=2.692 $X2=0
+ $Y2=0
cc_903 N_A_1355_377#_c_1355_n N_VPWR_c_1665_n 0.00851838f $X=7.01 $Y=2.692 $X2=0
+ $Y2=0
cc_904 N_A_1355_377#_c_1362_n N_VPWR_c_1665_n 0.00626376f $X=7.73 $Y=2.35 $X2=0
+ $Y2=0
cc_905 N_A_1355_377#_c_1348_n N_VPWR_c_1671_n 0.00461464f $X=9.475 $Y=2.465
+ $X2=0 $Y2=0
cc_906 N_A_1355_377#_c_1357_n N_VPWR_c_1671_n 0.0145938f $X=8.605 $Y=2.75 $X2=0
+ $Y2=0
cc_907 N_A_1355_377#_c_1349_n N_VPWR_c_1672_n 0.00444681f $X=9.98 $Y=1.765 $X2=0
+ $Y2=0
cc_908 N_A_1355_377#_c_1352_n N_VPWR_c_1672_n 0.00452264f $X=10.99 $Y=1.94 $X2=0
+ $Y2=0
cc_909 N_A_1355_377#_c_1348_n N_VPWR_c_1657_n 0.00450799f $X=9.475 $Y=2.465
+ $X2=0 $Y2=0
cc_910 N_A_1355_377#_c_1349_n N_VPWR_c_1657_n 0.00882517f $X=9.98 $Y=1.765 $X2=0
+ $Y2=0
cc_911 N_A_1355_377#_c_1352_n N_VPWR_c_1657_n 0.00465044f $X=10.99 $Y=1.94 $X2=0
+ $Y2=0
cc_912 N_A_1355_377#_c_1354_n N_VPWR_c_1657_n 0.0151143f $X=7.238 $Y=2.692 $X2=0
+ $Y2=0
cc_913 N_A_1355_377#_c_1355_n N_VPWR_c_1657_n 0.00866988f $X=7.01 $Y=2.692 $X2=0
+ $Y2=0
cc_914 N_A_1355_377#_c_1356_n N_VPWR_c_1657_n 0.0126283f $X=8.44 $Y=2.265 $X2=0
+ $Y2=0
cc_915 N_A_1355_377#_c_1357_n N_VPWR_c_1657_n 0.0120466f $X=8.605 $Y=2.75 $X2=0
+ $Y2=0
cc_916 N_A_1355_377#_c_1362_n N_VPWR_c_1657_n 0.0117647f $X=7.73 $Y=2.35 $X2=0
+ $Y2=0
cc_917 N_A_1355_377#_c_1362_n A_1517_508# 0.00159274f $X=7.73 $Y=2.35 $X2=-0.19
+ $Y2=-0.245
cc_918 N_A_1355_377#_c_1363_n A_1517_508# 0.00130139f $X=7.9 $Y=2.35 $X2=-0.19
+ $Y2=-0.245
cc_919 N_A_1355_377#_c_1337_n N_Q_N_c_1803_n 0.0141919f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_920 N_A_1355_377#_M1026_g N_Q_N_c_1803_n 0.00158934f $X=10.925 $Y=0.645 $X2=0
+ $Y2=0
cc_921 N_A_1355_377#_c_1349_n Q_N 0.0126086f $X=9.98 $Y=1.765 $X2=0 $Y2=0
cc_922 N_A_1355_377#_c_1338_n Q_N 0.0263745f $X=10.85 $Y=1.41 $X2=0 $Y2=0
cc_923 N_A_1355_377#_c_1339_n Q_N 0.00414194f $X=10.07 $Y=1.41 $X2=0 $Y2=0
cc_924 N_A_1355_377#_c_1352_n Q_N 0.00362081f $X=10.99 $Y=1.94 $X2=0 $Y2=0
cc_925 N_A_1355_377#_c_1337_n N_Q_N_c_1805_n 0.00565895f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_926 N_A_1355_377#_c_1338_n N_Q_N_c_1805_n 0.016272f $X=10.85 $Y=1.41 $X2=0
+ $Y2=0
cc_927 N_A_1355_377#_M1026_g N_Q_N_c_1805_n 0.00117107f $X=10.925 $Y=0.645 $X2=0
+ $Y2=0
cc_928 N_A_1355_377#_M1026_g N_Q_c_1834_n 6.13748e-19 $X=10.925 $Y=0.645 $X2=0
+ $Y2=0
cc_929 N_A_1355_377#_c_1352_n Q 6.18336e-19 $X=10.99 $Y=1.94 $X2=0 $Y2=0
cc_930 N_A_1355_377#_c_1353_n Q 5.87905e-19 $X=10.99 $Y=1.865 $X2=0 $Y2=0
cc_931 N_A_1355_377#_c_1334_n N_VGND_c_1859_n 0.00403474f $X=8.875 $Y=0.865
+ $X2=0 $Y2=0
cc_932 N_A_1355_377#_c_1337_n N_VGND_c_1859_n 0.0109009f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_933 N_A_1355_377#_c_1339_n N_VGND_c_1859_n 0.00184725f $X=10.07 $Y=1.41 $X2=0
+ $Y2=0
cc_934 N_A_1355_377#_M1026_g N_VGND_c_1860_n 0.00686847f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_935 N_A_1355_377#_c_1334_n N_VGND_c_1863_n 0.00435647f $X=8.875 $Y=0.865
+ $X2=0 $Y2=0
cc_936 N_A_1355_377#_c_1337_n N_VGND_c_1868_n 0.00434272f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_937 N_A_1355_377#_M1026_g N_VGND_c_1868_n 0.00434272f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_938 N_A_1355_377#_c_1334_n N_VGND_c_1870_n 0.00454088f $X=8.875 $Y=0.865
+ $X2=0 $Y2=0
cc_939 N_A_1355_377#_c_1337_n N_VGND_c_1870_n 0.00830058f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_940 N_A_1355_377#_M1026_g N_VGND_c_1870_n 0.00826607f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_941 N_A_1355_377#_c_1334_n N_VGND_c_1874_n 0.0074138f $X=8.875 $Y=0.865 $X2=0
+ $Y2=0
cc_942 N_A_2113_74#_c_1534_n N_VPWR_c_1664_n 0.0122635f $X=11.495 $Y=1.765 $X2=0
+ $Y2=0
cc_943 N_A_2113_74#_c_1538_n N_VPWR_c_1664_n 0.0573751f $X=10.765 $Y=2.16 $X2=0
+ $Y2=0
cc_944 N_A_2113_74#_c_1539_n N_VPWR_c_1664_n 0.0135101f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_945 N_A_2113_74#_c_1538_n N_VPWR_c_1672_n 0.00525601f $X=10.765 $Y=2.16 $X2=0
+ $Y2=0
cc_946 N_A_2113_74#_c_1534_n N_VPWR_c_1673_n 0.00445602f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_947 N_A_2113_74#_c_1534_n N_VPWR_c_1657_n 0.00865325f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_948 N_A_2113_74#_c_1538_n N_VPWR_c_1657_n 0.00579841f $X=10.765 $Y=2.16 $X2=0
+ $Y2=0
cc_949 N_A_2113_74#_c_1536_n N_Q_N_c_1803_n 0.0397432f $X=10.71 $Y=0.645 $X2=0
+ $Y2=0
cc_950 N_A_2113_74#_c_1537_n N_Q_N_c_1803_n 0.00113323f $X=10.777 $Y=1.22 $X2=0
+ $Y2=0
cc_951 N_A_2113_74#_c_1538_n Q_N 0.0793992f $X=10.765 $Y=2.16 $X2=0 $Y2=0
cc_952 N_A_2113_74#_c_1560_n Q_N 0.0126081f $X=10.777 $Y=1.385 $X2=0 $Y2=0
cc_953 N_A_2113_74#_c_1537_n N_Q_N_c_1805_n 0.0124563f $X=10.777 $Y=1.22 $X2=0
+ $Y2=0
cc_954 N_A_2113_74#_c_1560_n N_Q_N_c_1805_n 0.00696689f $X=10.777 $Y=1.385 $X2=0
+ $Y2=0
cc_955 N_A_2113_74#_c_1535_n N_Q_c_1834_n 0.00613596f $X=11.505 $Y=1.22 $X2=0
+ $Y2=0
cc_956 N_A_2113_74#_c_1535_n N_Q_c_1835_n 0.00402186f $X=11.505 $Y=1.22 $X2=0
+ $Y2=0
cc_957 N_A_2113_74#_c_1534_n Q 0.0162052f $X=11.495 $Y=1.765 $X2=0 $Y2=0
cc_958 N_A_2113_74#_c_1534_n N_Q_c_1836_n 0.0158104f $X=11.495 $Y=1.765 $X2=0
+ $Y2=0
cc_959 N_A_2113_74#_c_1535_n N_Q_c_1836_n 0.00424967f $X=11.505 $Y=1.22 $X2=0
+ $Y2=0
cc_960 N_A_2113_74#_c_1539_n N_Q_c_1836_n 0.0256386f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_961 N_A_2113_74#_c_1534_n N_VGND_c_1860_n 0.00278132f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_962 N_A_2113_74#_c_1535_n N_VGND_c_1860_n 0.00691628f $X=11.505 $Y=1.22 $X2=0
+ $Y2=0
cc_963 N_A_2113_74#_c_1536_n N_VGND_c_1860_n 0.022629f $X=10.71 $Y=0.645 $X2=0
+ $Y2=0
cc_964 N_A_2113_74#_c_1539_n N_VGND_c_1860_n 0.0190052f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_965 N_A_2113_74#_c_1536_n N_VGND_c_1868_n 0.0145025f $X=10.71 $Y=0.645 $X2=0
+ $Y2=0
cc_966 N_A_2113_74#_c_1535_n N_VGND_c_1869_n 0.00434272f $X=11.505 $Y=1.22 $X2=0
+ $Y2=0
cc_967 N_A_2113_74#_c_1535_n N_VGND_c_1870_n 0.00825042f $X=11.505 $Y=1.22 $X2=0
+ $Y2=0
cc_968 N_A_2113_74#_c_1536_n N_VGND_c_1870_n 0.0119747f $X=10.71 $Y=0.645 $X2=0
+ $Y2=0
cc_969 N_A_27_80#_c_1597_n N_VPWR_M1027_d 0.00134035f $X=2.525 $Y=2.145 $X2=0
+ $Y2=0
cc_970 N_A_27_80#_c_1641_n N_VPWR_M1027_d 0.005034f $X=1.71 $Y=2.145 $X2=0 $Y2=0
cc_971 N_A_27_80#_c_1595_n N_VPWR_c_1658_n 0.0261795f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_972 N_A_27_80#_c_1596_n N_VPWR_c_1658_n 0.0195982f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_973 N_A_27_80#_c_1596_n N_VPWR_c_1659_n 0.00102433f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_974 N_A_27_80#_c_1597_n N_VPWR_c_1659_n 0.00268134f $X=2.525 $Y=2.145 $X2=0
+ $Y2=0
cc_975 N_A_27_80#_c_1641_n N_VPWR_c_1659_n 0.0124964f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_976 N_A_27_80#_c_1595_n N_VPWR_c_1667_n 0.011066f $X=0.28 $Y=2.75 $X2=0 $Y2=0
cc_977 N_A_27_80#_c_1595_n N_VPWR_c_1657_n 0.00915947f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_978 N_A_27_80#_c_1589_n N_VGND_c_1854_n 0.0172562f $X=0.28 $Y=0.61 $X2=0
+ $Y2=0
cc_979 N_A_27_80#_c_1589_n N_VGND_c_1865_n 0.00978756f $X=0.28 $Y=0.61 $X2=0
+ $Y2=0
cc_980 N_A_27_80#_c_1589_n N_VGND_c_1870_n 0.00895297f $X=0.28 $Y=0.61 $X2=0
+ $Y2=0
cc_981 N_VPWR_c_1663_n Q_N 0.0165387f $X=9.735 $Y=2.815 $X2=0 $Y2=0
cc_982 N_VPWR_c_1664_n Q_N 0.00312692f $X=11.215 $Y=2.16 $X2=0 $Y2=0
cc_983 N_VPWR_c_1672_n Q_N 0.0139663f $X=11.05 $Y=3.33 $X2=0 $Y2=0
cc_984 N_VPWR_c_1657_n Q_N 0.0115601f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_985 N_VPWR_c_1664_n Q 0.0368843f $X=11.215 $Y=2.16 $X2=0 $Y2=0
cc_986 N_VPWR_c_1673_n Q 0.0145938f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_987 N_VPWR_c_1657_n Q 0.0120466f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_988 N_Q_N_c_1803_n N_VGND_c_1859_n 0.0127977f $X=10.15 $Y=0.515 $X2=0 $Y2=0
cc_989 N_Q_N_c_1803_n N_VGND_c_1868_n 0.0145639f $X=10.15 $Y=0.515 $X2=0 $Y2=0
cc_990 N_Q_N_c_1803_n N_VGND_c_1870_n 0.0119984f $X=10.15 $Y=0.515 $X2=0 $Y2=0
cc_991 N_Q_c_1834_n N_VGND_c_1860_n 0.0228912f $X=11.72 $Y=0.515 $X2=0 $Y2=0
cc_992 N_Q_c_1834_n N_VGND_c_1869_n 0.0145787f $X=11.72 $Y=0.515 $X2=0 $Y2=0
cc_993 N_Q_c_1834_n N_VGND_c_1870_n 0.0120042f $X=11.72 $Y=0.515 $X2=0 $Y2=0
