* NGSPICE file created from sky130_fd_sc_hs__sedfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 a_661_113# a_631_87# a_1071_455# VPB pshort w=640000u l=150000u
+  ad=4.707e+11p pd=5.06e+06u as=1.536e+11p ps=1.76e+06u
M1001 VPWR DE a_177_290# VPB pshort w=640000u l=150000u
+  ad=3.30785e+12p pd=2.82e+07u as=1.888e+11p ps=1.87e+06u
M1002 a_135_74# D a_37_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.373e+11p ps=2.81e+06u
M1003 a_661_113# SCE a_1044_125# VNB nlowvt w=420000u l=150000u
+  ad=5.502e+11p pd=5.14e+06u as=8.82e+10p ps=1.26e+06u
M1004 VPWR a_2403_74# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1005 a_1756_97# a_1510_74# a_661_113# VPB pshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1006 a_2403_74# a_1313_74# a_2292_392# VPB pshort w=1e+06u l=150000u
+  ad=3.049e+11p pd=2.72e+06u as=8.1e+11p ps=3.62e+06u
M1007 VPWR a_1943_53# a_1899_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1008 VGND DE a_177_290# VNB nlowvt w=420000u l=150000u
+  ad=2.3264e+12p pd=2.159e+07u as=1.197e+11p ps=1.41e+06u
M1009 Q a_2403_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1899_508# a_1313_74# a_1756_97# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1044_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_2403_74# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1510_74# a_1313_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1014 a_2586_508# a_1510_74# a_2403_74# VPB pshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1015 a_37_464# a_545_87# a_572_463# VPB pshort w=640000u l=150000u
+  ad=3.808e+11p pd=3.75e+06u as=1.536e+11p ps=1.76e+06u
M1016 a_2498_74# a_1313_74# a_2403_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.915e+11p ps=1.93e+06u
M1017 VGND a_545_87# a_2498_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_126_464# D a_37_464# VPB pshort w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1019 a_661_113# SCE a_37_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_545_87# a_2403_74# VPWR VPB pshort w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=0p ps=0u
M1021 a_545_87# a_2403_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1022 Q a_2403_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.255e+11p pd=4.11e+06u as=0p ps=0u
M1023 a_37_464# a_545_87# a_497_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1024 a_661_113# a_631_87# a_37_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1313_74# CLK VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1026 a_1313_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1027 a_2292_392# a_1943_53# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Q a_2403_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1510_74# a_1313_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1030 a_572_463# DE VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2403_74# a_1510_74# a_2331_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1032 VGND a_1943_53# a_1858_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.785e+11p ps=1.69e+06u
M1033 a_1071_455# SCD VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND DE a_135_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_545_87# a_2586_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1858_79# a_1510_74# a_1756_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.6695e+11p ps=1.74e+06u
M1037 VPWR a_177_290# a_126_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_497_113# a_177_290# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_2403_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1756_97# a_1313_74# a_661_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_2403_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 Q a_2403_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1943_53# a_1756_97# VPWR VPB pshort w=840000u l=150000u
+  ad=2.31e+11p pd=2.23e+06u as=0p ps=0u
M1044 VPWR SCE a_631_87# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1045 VGND SCE a_631_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1046 a_1943_53# a_1756_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1047 a_2331_74# a_1943_53# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

