* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 a_1278_121# a_758_306# a_1191_121# VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=9.2755e+11p ps=8.21e+06u
M1001 a_1191_121# a_758_306# a_1278_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_509_392# S0 a_114_126# VNB nlowvt w=640000u l=150000u
+  ad=8.5705e+11p pd=8.11e+06u as=3.872e+11p ps=3.77e+06u
M1003 VPWR S1 a_2489_347# VPB pshort w=1.12e+06u l=150000u
+  ad=3.70125e+12p pd=2.87e+07u as=3.696e+11p ps=2.9e+06u
M1004 a_1450_121# S0 a_1191_121# VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1005 a_1285_377# a_758_306# a_1191_121# VPB pshort w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=1.24e+12p ps=1.048e+07u
M1006 VPWR A3 a_1285_377# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_2199_74# a_2489_347# a_1191_121# VPB pshort w=1e+06u l=150000u
+  ad=9.9e+11p pd=7.98e+06u as=0p ps=0u
M1008 a_1191_121# a_758_306# a_1285_377# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1191_121# a_2489_347# a_2199_74# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND S1 a_2489_347# VNB nlowvt w=740000u l=150000u
+  ad=2.4642e+12p pd=2.151e+07u as=2.109e+11p ps=2.05e+06u
M1011 a_509_392# S1 a_2199_74# VPB pshort w=1e+06u l=150000u
+  ad=1.28e+12p pd=1.056e+07u as=0p ps=0u
M1012 a_2199_74# S1 a_509_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_2199_74# a_2489_347# a_509_392# VNB nlowvt w=640000u l=150000u
+  ad=8.576e+11p pd=6.52e+06u as=0p ps=0u
M1014 a_1465_377# S0 a_1191_121# VPB pshort w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1015 a_116_392# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1016 VPWR A1 a_116_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_509_392# S0 a_296_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=6.75e+11p ps=5.35e+06u
M1018 VGND S0 a_758_306# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1019 X a_2199_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1020 a_1191_121# S1 a_2199_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_296_392# A0 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A0 a_296_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1191_121# S0 a_1465_377# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1450_121# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2199_74# S1 a_1191_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_2199_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1027 a_1278_121# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_296_392# S0 a_509_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR S0 a_758_306# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1030 a_299_126# A0 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1031 a_116_392# a_758_306# a_509_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND A0 a_299_126# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_509_392# a_758_306# a_116_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A1 a_114_126# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_2199_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND A3 a_1450_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_114_126# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_2199_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1285_377# A3 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_299_126# a_758_306# a_509_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND A2 a_1278_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1191_121# S0 a_1450_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 X a_2199_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_509_392# a_758_306# a_299_126# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR a_2199_74# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1465_377# A2 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_114_126# S0 a_509_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 VPWR a_2199_74# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_509_392# a_2489_347# a_2199_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VPWR A2 a_1465_377# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 X a_2199_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
