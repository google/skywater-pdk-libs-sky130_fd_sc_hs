* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 Q a_821_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_1449_368# a_821_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_569_80# a_363_82# a_641_80# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 Q a_821_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR a_27_112# a_566_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_821_98# a_641_80# a_1049_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND a_821_98# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR a_641_80# a_821_98# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 a_641_80# a_230_74# a_773_124# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 VPWR GATE a_230_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 a_641_80# a_363_82# a_757_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 a_27_112# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X12 a_757_508# a_821_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X13 a_363_82# a_230_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_821_98# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X15 VGND a_27_112# a_569_80# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 VGND a_1449_368# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VPWR a_821_98# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X18 Q_N a_1449_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X19 a_1449_368# a_821_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_27_112# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X21 VGND GATE a_230_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 Q_N a_1449_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_1049_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_566_392# a_230_74# a_641_80# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X25 a_773_124# a_821_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 VPWR a_1449_368# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X27 a_363_82# a_230_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
.ends
