* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_376_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 VPWR B1 a_376_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 a_776_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 a_311_85# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 Y C1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_311_85# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_27_74# B1 a_311_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_27_74# B2 a_311_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_311_85# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VGND A2 a_311_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 Y A2 a_776_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X12 a_311_85# B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X14 a_776_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X15 Y B2 a_376_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 a_376_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X17 VPWR A1 a_776_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X18 a_27_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VGND A1 a_311_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
