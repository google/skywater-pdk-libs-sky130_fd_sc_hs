* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_83_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 VPWR A1 a_346_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_83_264# B2 a_652_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 a_83_264# B1 a_349_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_652_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 VGND A1 a_349_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_430_368# A3 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X8 a_349_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X10 a_349_74# B2 a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_346_368# A2 a_430_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X12 VGND a_83_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VGND A3 a_349_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
