* File: sky130_fd_sc_hs__a21o_2.pxi.spice
* Created: Tue Sep  1 19:49:39 2020
* 
x_PM_SKY130_FD_SC_HS__A21O_2%A_84_244# N_A_84_244#_M1004_d N_A_84_244#_M1003_s
+ N_A_84_244#_c_67_n N_A_84_244#_M1001_g N_A_84_244#_c_60_n N_A_84_244#_M1000_g
+ N_A_84_244#_c_68_n N_A_84_244#_M1002_g N_A_84_244#_c_61_n N_A_84_244#_M1007_g
+ N_A_84_244#_c_62_n N_A_84_244#_c_63_n N_A_84_244#_c_77_p N_A_84_244#_c_128_p
+ N_A_84_244#_c_70_n N_A_84_244#_c_71_n N_A_84_244#_c_64_n N_A_84_244#_c_65_n
+ N_A_84_244#_c_66_n PM_SKY130_FD_SC_HS__A21O_2%A_84_244#
x_PM_SKY130_FD_SC_HS__A21O_2%B1 N_B1_M1004_g N_B1_M1003_g N_B1_c_147_n
+ N_B1_c_152_n B1 N_B1_c_148_n N_B1_c_149_n N_B1_c_150_n
+ PM_SKY130_FD_SC_HS__A21O_2%B1
x_PM_SKY130_FD_SC_HS__A21O_2%A1 N_A1_M1009_g N_A1_c_186_n N_A1_c_191_n
+ N_A1_M1005_g A1 N_A1_c_188_n N_A1_c_189_n PM_SKY130_FD_SC_HS__A21O_2%A1
x_PM_SKY130_FD_SC_HS__A21O_2%A2 N_A2_c_226_n N_A2_M1008_g N_A2_M1006_g
+ N_A2_c_227_n N_A2_c_231_n A2 N_A2_c_229_n PM_SKY130_FD_SC_HS__A21O_2%A2
x_PM_SKY130_FD_SC_HS__A21O_2%VPWR N_VPWR_M1001_d N_VPWR_M1002_d N_VPWR_M1005_d
+ N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n N_VPWR_c_260_n VPWR
+ N_VPWR_c_261_n N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_256_n N_VPWR_c_265_n
+ N_VPWR_c_266_n PM_SKY130_FD_SC_HS__A21O_2%VPWR
x_PM_SKY130_FD_SC_HS__A21O_2%X N_X_M1000_d N_X_M1001_s N_X_c_300_n N_X_c_305_n X
+ X X X N_X_c_301_n PM_SKY130_FD_SC_HS__A21O_2%X
x_PM_SKY130_FD_SC_HS__A21O_2%A_401_392# N_A_401_392#_M1003_d
+ N_A_401_392#_M1006_d N_A_401_392#_c_329_n N_A_401_392#_c_330_n
+ N_A_401_392#_c_331_n N_A_401_392#_c_332_n
+ PM_SKY130_FD_SC_HS__A21O_2%A_401_392#
x_PM_SKY130_FD_SC_HS__A21O_2%VGND N_VGND_M1000_s N_VGND_M1007_s N_VGND_M1008_d
+ N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n
+ N_VGND_c_363_n VGND N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n
+ N_VGND_c_367_n PM_SKY130_FD_SC_HS__A21O_2%VGND
cc_1 VNB N_A_84_244#_c_60_n 0.0199304f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.22
cc_2 VNB N_A_84_244#_c_61_n 0.0197587f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.22
cc_3 VNB N_A_84_244#_c_62_n 0.00175887f $X=-0.19 $Y=-0.245 $X2=1.232 $Y2=1.382
cc_4 VNB N_A_84_244#_c_63_n 0.00209425f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.385
cc_5 VNB N_A_84_244#_c_64_n 0.0024006f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=0.495
cc_6 VNB N_A_84_244#_c_65_n 0.00190688f $X=-0.19 $Y=-0.245 $X2=1.232 $Y2=1.22
cc_7 VNB N_A_84_244#_c_66_n 0.100903f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.492
cc_8 VNB N_B1_c_147_n 0.00686523f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_9 VNB N_B1_c_148_n 0.0300812f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_10 VNB N_B1_c_149_n 0.00796318f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_11 VNB N_B1_c_150_n 0.0198297f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.22
cc_12 VNB N_A1_c_186_n 0.0064486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A1 0.0172207f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_14 VNB N_A1_c_188_n 0.0270606f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.74
cc_15 VNB N_A1_c_189_n 0.0177861f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_16 VNB N_A2_c_226_n 0.0212479f $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=0.37
cc_17 VNB N_A2_c_227_n 0.00903934f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_18 VNB A2 0.0104864f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.74
cc_19 VNB N_A2_c_229_n 0.0594649f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.74
cc_20 VNB N_VPWR_c_256_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.492
cc_21 VNB N_X_c_300_n 0.00240251f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_22 VNB N_X_c_301_n 8.09729e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_358_n 0.0474446f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.74
cc_24 VNB N_VGND_c_359_n 0.0123902f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.22
cc_25 VNB N_VGND_c_360_n 0.0136221f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.74
cc_26 VNB N_VGND_c_361_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=1.232 $Y2=1.705
cc_27 VNB N_VGND_c_362_n 0.0115308f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.385
cc_28 VNB N_VGND_c_363_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.01
cc_29 VNB N_VGND_c_364_n 0.019013f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=2.105
cc_30 VNB N_VGND_c_365_n 0.0312656f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=0.84
cc_31 VNB N_VGND_c_366_n 0.0109638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_367_n 0.22003f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.492
cc_33 VPB N_A_84_244#_c_67_n 0.0174317f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_34 VPB N_A_84_244#_c_68_n 0.0168737f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_35 VPB N_A_84_244#_c_63_n 0.00177895f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.385
cc_36 VPB N_A_84_244#_c_70_n 0.0213178f $X=-0.19 $Y=1.66 $X2=1.665 $Y2=1.875
cc_37 VPB N_A_84_244#_c_71_n 0.0150325f $X=-0.19 $Y=1.66 $X2=1.705 $Y2=2.105
cc_38 VPB N_A_84_244#_c_66_n 0.0160637f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=1.492
cc_39 VPB N_B1_c_147_n 0.00721108f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_40 VPB N_B1_c_152_n 0.0231102f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.22
cc_41 VPB N_A1_c_186_n 0.00695588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A1_c_191_n 0.0203815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A2_c_227_n 0.00905166f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_44 VPB N_A2_c_231_n 0.0247613f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.22
cc_45 VPB N_VPWR_c_257_n 0.0108116f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.22
cc_46 VPB N_VPWR_c_258_n 0.0647053f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=0.74
cc_47 VPB N_VPWR_c_259_n 0.0149716f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=0.74
cc_48 VPB N_VPWR_c_260_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.01
cc_49 VPB N_VPWR_c_261_n 0.0182909f $X=-0.19 $Y=1.66 $X2=1.705 $Y2=2.105
cc_50 VPB N_VPWR_c_262_n 0.0305896f $X=-0.19 $Y=1.66 $X2=2.13 $Y2=0.495
cc_51 VPB N_VPWR_c_263_n 0.0188229f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_256_n 0.074034f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.492
cc_53 VPB N_VPWR_c_265_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_266_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB X 0.00243101f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_56 VPB N_A_401_392#_c_329_n 0.00282887f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_57 VPB N_A_401_392#_c_330_n 0.0194475f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_58 VPB N_A_401_392#_c_331_n 0.00879836f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_59 VPB N_A_401_392#_c_332_n 0.0440661f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=0.74
cc_60 N_A_84_244#_c_63_n N_B1_c_147_n 0.004282f $X=1.23 $Y=1.385 $X2=0 $Y2=0
cc_61 N_A_84_244#_c_70_n N_B1_c_147_n 0.00433566f $X=1.665 $Y=1.875 $X2=0 $Y2=0
cc_62 N_A_84_244#_c_71_n N_B1_c_152_n 0.00578804f $X=1.705 $Y=2.105 $X2=0 $Y2=0
cc_63 N_A_84_244#_c_62_n N_B1_c_148_n 3.35236e-19 $X=1.232 $Y=1.382 $X2=0 $Y2=0
cc_64 N_A_84_244#_c_77_p N_B1_c_148_n 0.00102115f $X=1.965 $Y=0.925 $X2=0 $Y2=0
cc_65 N_A_84_244#_c_70_n N_B1_c_148_n 0.00296638f $X=1.665 $Y=1.875 $X2=0 $Y2=0
cc_66 N_A_84_244#_c_66_n N_B1_c_148_n 0.0163108f $X=1.105 $Y=1.492 $X2=0 $Y2=0
cc_67 N_A_84_244#_c_77_p N_B1_c_149_n 0.0303988f $X=1.965 $Y=0.925 $X2=0 $Y2=0
cc_68 N_A_84_244#_c_70_n N_B1_c_149_n 0.017401f $X=1.665 $Y=1.875 $X2=0 $Y2=0
cc_69 N_A_84_244#_c_65_n N_B1_c_149_n 0.0285482f $X=1.232 $Y=1.22 $X2=0 $Y2=0
cc_70 N_A_84_244#_c_66_n N_B1_c_149_n 0.00227878f $X=1.105 $Y=1.492 $X2=0 $Y2=0
cc_71 N_A_84_244#_c_61_n N_B1_c_150_n 0.00826871f $X=1.105 $Y=1.22 $X2=0 $Y2=0
cc_72 N_A_84_244#_c_77_p N_B1_c_150_n 0.0105649f $X=1.965 $Y=0.925 $X2=0 $Y2=0
cc_73 N_A_84_244#_c_64_n N_B1_c_150_n 0.0116638f $X=2.13 $Y=0.495 $X2=0 $Y2=0
cc_74 N_A_84_244#_c_65_n N_B1_c_150_n 0.00301427f $X=1.232 $Y=1.22 $X2=0 $Y2=0
cc_75 N_A_84_244#_c_77_p A1 0.00552432f $X=1.965 $Y=0.925 $X2=0 $Y2=0
cc_76 N_A_84_244#_c_77_p N_A1_c_188_n 3.3691e-19 $X=1.965 $Y=0.925 $X2=0 $Y2=0
cc_77 N_A_84_244#_c_77_p N_A1_c_189_n 0.00339533f $X=1.965 $Y=0.925 $X2=0 $Y2=0
cc_78 N_A_84_244#_c_64_n N_A1_c_189_n 0.00988058f $X=2.13 $Y=0.495 $X2=0 $Y2=0
cc_79 N_A_84_244#_c_77_p N_A2_c_226_n 5.12803e-19 $X=1.965 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_84_244#_c_64_n N_A2_c_226_n 0.00148221f $X=2.13 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_81 N_A_84_244#_c_70_n N_VPWR_M1002_d 0.00266686f $X=1.665 $Y=1.875 $X2=0
+ $Y2=0
cc_82 N_A_84_244#_c_67_n N_VPWR_c_258_n 0.008783f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_84_244#_c_67_n N_VPWR_c_259_n 6.11953e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_84_244#_c_68_n N_VPWR_c_259_n 0.0144702f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_84_244#_c_70_n N_VPWR_c_259_n 0.0210301f $X=1.665 $Y=1.875 $X2=0 $Y2=0
cc_86 N_A_84_244#_c_71_n N_VPWR_c_259_n 0.0705155f $X=1.705 $Y=2.105 $X2=0 $Y2=0
cc_87 N_A_84_244#_c_67_n N_VPWR_c_261_n 0.00445602f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_84_244#_c_68_n N_VPWR_c_261_n 0.00413917f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_84_244#_c_71_n N_VPWR_c_262_n 0.011066f $X=1.705 $Y=2.105 $X2=0 $Y2=0
cc_90 N_A_84_244#_c_67_n N_VPWR_c_256_n 0.008611f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_84_244#_c_68_n N_VPWR_c_256_n 0.00817726f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_84_244#_c_71_n N_VPWR_c_256_n 0.00915947f $X=1.705 $Y=2.105 $X2=0
+ $Y2=0
cc_93 N_A_84_244#_c_60_n N_X_c_300_n 0.00629186f $X=0.675 $Y=1.22 $X2=0 $Y2=0
cc_94 N_A_84_244#_c_61_n N_X_c_300_n 0.0117096f $X=1.105 $Y=1.22 $X2=0 $Y2=0
cc_95 N_A_84_244#_c_60_n N_X_c_305_n 0.00180034f $X=0.675 $Y=1.22 $X2=0 $Y2=0
cc_96 N_A_84_244#_c_61_n N_X_c_305_n 0.00295249f $X=1.105 $Y=1.22 $X2=0 $Y2=0
cc_97 N_A_84_244#_c_66_n N_X_c_305_n 0.00192922f $X=1.105 $Y=1.492 $X2=0 $Y2=0
cc_98 N_A_84_244#_c_67_n X 0.00397951f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_84_244#_c_68_n X 0.00299619f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_84_244#_c_63_n X 0.0178828f $X=1.23 $Y=1.385 $X2=0 $Y2=0
cc_101 N_A_84_244#_c_70_n X 0.0125498f $X=1.665 $Y=1.875 $X2=0 $Y2=0
cc_102 N_A_84_244#_c_71_n X 4.23899e-19 $X=1.705 $Y=2.105 $X2=0 $Y2=0
cc_103 N_A_84_244#_c_66_n X 0.0277563f $X=1.105 $Y=1.492 $X2=0 $Y2=0
cc_104 N_A_84_244#_c_67_n X 0.0125514f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_84_244#_c_68_n X 3.88029e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A_84_244#_c_60_n N_X_c_301_n 0.0054987f $X=0.675 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A_84_244#_c_61_n N_X_c_301_n 0.00122577f $X=1.105 $Y=1.22 $X2=0 $Y2=0
cc_108 N_A_84_244#_c_62_n N_X_c_301_n 0.0178828f $X=1.232 $Y=1.382 $X2=0 $Y2=0
cc_109 N_A_84_244#_c_65_n N_X_c_301_n 0.00657203f $X=1.232 $Y=1.22 $X2=0 $Y2=0
cc_110 N_A_84_244#_c_66_n N_X_c_301_n 0.0245841f $X=1.105 $Y=1.492 $X2=0 $Y2=0
cc_111 N_A_84_244#_c_71_n N_A_401_392#_c_329_n 0.0716912f $X=1.705 $Y=2.105
+ $X2=0 $Y2=0
cc_112 N_A_84_244#_c_70_n N_A_401_392#_c_331_n 0.0121546f $X=1.665 $Y=1.875
+ $X2=0 $Y2=0
cc_113 N_A_84_244#_c_71_n N_A_401_392#_c_331_n 0.00105301f $X=1.705 $Y=2.105
+ $X2=0 $Y2=0
cc_114 N_A_84_244#_c_77_p N_VGND_M1007_s 0.0150178f $X=1.965 $Y=0.925 $X2=0
+ $Y2=0
cc_115 N_A_84_244#_c_128_p N_VGND_M1007_s 0.00321143f $X=1.395 $Y=0.925 $X2=0
+ $Y2=0
cc_116 N_A_84_244#_c_65_n N_VGND_M1007_s 0.00170409f $X=1.232 $Y=1.22 $X2=0
+ $Y2=0
cc_117 N_A_84_244#_c_60_n N_VGND_c_358_n 0.00647412f $X=0.675 $Y=1.22 $X2=0
+ $Y2=0
cc_118 N_A_84_244#_c_66_n N_VGND_c_358_n 0.00652095f $X=1.105 $Y=1.492 $X2=0
+ $Y2=0
cc_119 N_A_84_244#_c_61_n N_VGND_c_359_n 0.00404337f $X=1.105 $Y=1.22 $X2=0
+ $Y2=0
cc_120 N_A_84_244#_c_77_p N_VGND_c_359_n 0.0308408f $X=1.965 $Y=0.925 $X2=0
+ $Y2=0
cc_121 N_A_84_244#_c_128_p N_VGND_c_359_n 0.0139023f $X=1.395 $Y=0.925 $X2=0
+ $Y2=0
cc_122 N_A_84_244#_c_64_n N_VGND_c_359_n 0.0128657f $X=2.13 $Y=0.495 $X2=0 $Y2=0
cc_123 N_A_84_244#_c_66_n N_VGND_c_359_n 5.89585e-19 $X=1.105 $Y=1.492 $X2=0
+ $Y2=0
cc_124 N_A_84_244#_c_77_p N_VGND_c_361_n 0.00499344f $X=1.965 $Y=0.925 $X2=0
+ $Y2=0
cc_125 N_A_84_244#_c_64_n N_VGND_c_361_n 0.0135598f $X=2.13 $Y=0.495 $X2=0 $Y2=0
cc_126 N_A_84_244#_c_60_n N_VGND_c_364_n 0.00434272f $X=0.675 $Y=1.22 $X2=0
+ $Y2=0
cc_127 N_A_84_244#_c_61_n N_VGND_c_364_n 0.00434272f $X=1.105 $Y=1.22 $X2=0
+ $Y2=0
cc_128 N_A_84_244#_c_64_n N_VGND_c_365_n 0.0144609f $X=2.13 $Y=0.495 $X2=0 $Y2=0
cc_129 N_A_84_244#_c_60_n N_VGND_c_367_n 0.00824418f $X=0.675 $Y=1.22 $X2=0
+ $Y2=0
cc_130 N_A_84_244#_c_61_n N_VGND_c_367_n 0.0082272f $X=1.105 $Y=1.22 $X2=0 $Y2=0
cc_131 N_A_84_244#_c_77_p N_VGND_c_367_n 0.00627901f $X=1.965 $Y=0.925 $X2=0
+ $Y2=0
cc_132 N_A_84_244#_c_128_p N_VGND_c_367_n 6.15084e-19 $X=1.395 $Y=0.925 $X2=0
+ $Y2=0
cc_133 N_A_84_244#_c_64_n N_VGND_c_367_n 0.0118703f $X=2.13 $Y=0.495 $X2=0 $Y2=0
cc_134 N_B1_c_147_n N_A1_c_186_n 0.0109801f $X=1.922 $Y=1.79 $X2=0 $Y2=0
cc_135 N_B1_c_152_n N_A1_c_186_n 0.00416562f $X=1.922 $Y=1.885 $X2=0 $Y2=0
cc_136 N_B1_c_152_n N_A1_c_191_n 0.00815318f $X=1.922 $Y=1.885 $X2=0 $Y2=0
cc_137 N_B1_c_148_n A1 5.01118e-19 $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_138 N_B1_c_149_n A1 0.0240773f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_139 N_B1_c_148_n N_A1_c_188_n 0.0213922f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_140 N_B1_c_149_n N_A1_c_188_n 3.95971e-19 $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_141 N_B1_c_150_n N_A1_c_189_n 0.0131285f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_142 N_B1_c_152_n N_VPWR_c_259_n 0.00424964f $X=1.922 $Y=1.885 $X2=0 $Y2=0
cc_143 N_B1_c_152_n N_VPWR_c_260_n 8.23897e-19 $X=1.922 $Y=1.885 $X2=0 $Y2=0
cc_144 N_B1_c_152_n N_VPWR_c_262_n 0.00445602f $X=1.922 $Y=1.885 $X2=0 $Y2=0
cc_145 N_B1_c_152_n N_VPWR_c_256_n 0.00863237f $X=1.922 $Y=1.885 $X2=0 $Y2=0
cc_146 N_B1_c_152_n N_A_401_392#_c_329_n 0.0126899f $X=1.922 $Y=1.885 $X2=0
+ $Y2=0
cc_147 N_B1_c_147_n N_A_401_392#_c_331_n 6.92951e-19 $X=1.922 $Y=1.79 $X2=0
+ $Y2=0
cc_148 N_B1_c_152_n N_A_401_392#_c_331_n 0.00241612f $X=1.922 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_B1_c_150_n N_VGND_c_359_n 0.00404337f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_150 N_B1_c_150_n N_VGND_c_365_n 0.00434272f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_151 N_B1_c_150_n N_VGND_c_367_n 0.00447595f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_152 A1 N_A2_c_226_n 0.00160391f $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_153 N_A1_c_189_n N_A2_c_226_n 0.0363226f $X=2.365 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A1_c_186_n N_A2_c_227_n 0.0110538f $X=2.38 $Y=1.795 $X2=0 $Y2=0
cc_155 N_A1_c_186_n N_A2_c_231_n 0.00416562f $X=2.38 $Y=1.795 $X2=0 $Y2=0
cc_156 N_A1_c_191_n N_A2_c_231_n 0.00825045f $X=2.38 $Y=1.885 $X2=0 $Y2=0
cc_157 A1 A2 0.0290219f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A1_c_188_n A2 2.10483e-19 $X=2.365 $Y=1.385 $X2=0 $Y2=0
cc_159 A1 N_A2_c_229_n 0.00826783f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A1_c_188_n N_A2_c_229_n 0.0214735f $X=2.365 $Y=1.385 $X2=0 $Y2=0
cc_161 N_A1_c_191_n N_VPWR_c_260_n 0.0133917f $X=2.38 $Y=1.885 $X2=0 $Y2=0
cc_162 N_A1_c_191_n N_VPWR_c_262_n 0.00413917f $X=2.38 $Y=1.885 $X2=0 $Y2=0
cc_163 N_A1_c_191_n N_VPWR_c_256_n 0.0081781f $X=2.38 $Y=1.885 $X2=0 $Y2=0
cc_164 N_A1_c_191_n N_A_401_392#_c_329_n 0.00715681f $X=2.38 $Y=1.885 $X2=0
+ $Y2=0
cc_165 N_A1_c_186_n N_A_401_392#_c_330_n 0.00541098f $X=2.38 $Y=1.795 $X2=0
+ $Y2=0
cc_166 N_A1_c_191_n N_A_401_392#_c_330_n 0.0103148f $X=2.38 $Y=1.885 $X2=0 $Y2=0
cc_167 A1 N_A_401_392#_c_330_n 0.0392159f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_168 N_A1_c_188_n N_A_401_392#_c_330_n 0.00254286f $X=2.365 $Y=1.385 $X2=0
+ $Y2=0
cc_169 A1 N_A_401_392#_c_331_n 0.00339997f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A1_c_188_n N_A_401_392#_c_331_n 9.31826e-19 $X=2.365 $Y=1.385 $X2=0
+ $Y2=0
cc_171 N_A1_c_189_n N_VGND_c_361_n 0.00253696f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_172 N_A1_c_189_n N_VGND_c_365_n 0.00434272f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_173 N_A1_c_189_n N_VGND_c_367_n 0.00821825f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_174 N_A2_c_231_n N_VPWR_c_260_n 0.0165249f $X=2.837 $Y=1.885 $X2=0 $Y2=0
cc_175 N_A2_c_231_n N_VPWR_c_263_n 0.00413917f $X=2.837 $Y=1.885 $X2=0 $Y2=0
cc_176 N_A2_c_231_n N_VPWR_c_256_n 0.00821301f $X=2.837 $Y=1.885 $X2=0 $Y2=0
cc_177 N_A2_c_227_n N_A_401_392#_c_330_n 0.00972987f $X=2.837 $Y=1.79 $X2=0
+ $Y2=0
cc_178 N_A2_c_231_n N_A_401_392#_c_330_n 0.0110339f $X=2.837 $Y=1.885 $X2=0
+ $Y2=0
cc_179 A2 N_A_401_392#_c_330_n 0.0246672f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A2_c_229_n N_A_401_392#_c_330_n 0.00322993f $X=3.09 $Y=1.385 $X2=0
+ $Y2=0
cc_181 N_A2_c_231_n N_A_401_392#_c_332_n 0.00846769f $X=2.837 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_A2_c_226_n N_VGND_c_361_n 0.0188724f $X=2.815 $Y=1.22 $X2=0 $Y2=0
cc_183 A2 N_VGND_c_361_n 0.0226256f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A2_c_229_n N_VGND_c_361_n 0.00184416f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_185 N_A2_c_226_n N_VGND_c_365_n 0.00383152f $X=2.815 $Y=1.22 $X2=0 $Y2=0
cc_186 N_A2_c_226_n N_VGND_c_367_n 0.00757998f $X=2.815 $Y=1.22 $X2=0 $Y2=0
cc_187 N_VPWR_c_258_n X 0.0769137f $X=0.285 $Y=1.985 $X2=0 $Y2=0
cc_188 N_VPWR_c_259_n X 0.0358545f $X=1.185 $Y=2.13 $X2=0 $Y2=0
cc_189 N_VPWR_c_261_n X 0.0123628f $X=1.02 $Y=3.33 $X2=0 $Y2=0
cc_190 N_VPWR_c_256_n X 0.0101999f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_191 N_VPWR_c_260_n N_A_401_392#_c_329_n 0.0617165f $X=2.605 $Y=2.155 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_262_n N_A_401_392#_c_329_n 0.0110241f $X=2.44 $Y=3.33 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_256_n N_A_401_392#_c_329_n 0.00909194f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_260_n N_A_401_392#_c_330_n 0.021739f $X=2.605 $Y=2.155 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_260_n N_A_401_392#_c_332_n 0.0617165f $X=2.605 $Y=2.155 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_263_n N_A_401_392#_c_332_n 0.011066f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_256_n N_A_401_392#_c_332_n 0.00915947f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_198 N_X_c_300_n N_VGND_c_358_n 0.0290778f $X=0.89 $Y=0.515 $X2=0 $Y2=0
cc_199 N_X_c_300_n N_VGND_c_359_n 0.0128657f $X=0.89 $Y=0.515 $X2=0 $Y2=0
cc_200 N_X_c_300_n N_VGND_c_364_n 0.0145065f $X=0.89 $Y=0.515 $X2=0 $Y2=0
cc_201 N_X_c_300_n N_VGND_c_367_n 0.0118883f $X=0.89 $Y=0.515 $X2=0 $Y2=0
