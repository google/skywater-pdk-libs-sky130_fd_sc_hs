* File: sky130_fd_sc_hs__a222oi_1.spice
* Created: Tue Sep  1 19:50:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a222oi_1.pex.spice"
.subckt sky130_fd_sc_hs__a222oi_1  VNB VPB C1 C2 B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C2	C2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1007 A_119_74# N_C1_M1007_g N_Y_M1007_s VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2 SB=75003.5
+ A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_C2_M1000_g A_119_74# VNB NLOWVT L=0.15 W=0.64 AD=0.3744
+ AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75000.6 SB=75003.1
+ A=0.096 P=1.58 MULT=1
MM1005 A_461_74# N_B2_M1005_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.3744 PD=0.88 PS=1.81 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75001.9 SB=75001.8
+ A=0.096 P=1.58 MULT=1
MM1008 N_Y_M1008_d N_B1_M1008_g A_461_74# VNB NLOWVT L=0.15 W=0.64 AD=0.2048
+ AS=0.0768 PD=1.28 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75002.3 SB=75001.4
+ A=0.096 P=1.58 MULT=1
MM1010 A_697_74# N_A1_M1010_g N_Y_M1008_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.2048 PD=0.88 PS=1.28 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75003.1 SB=75000.6
+ A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g A_697_74# VNB NLOWVT L=0.15 W=0.64 AD=0.1824
+ AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75003.5 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1006 N_A_116_392#_M1006_d N_C1_M1006_g N_Y_M1006_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1003 N_Y_M1003_d N_C2_M1003_g N_A_116_392#_M1006_d VPB PSHORT L=0.15 W=1
+ AD=0.345 AS=0.175 PD=2.69 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1004 N_A_116_392#_M1004_d N_B2_M1004_g N_A_369_392#_M1004_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1001 N_A_369_392#_M1001_d N_B1_M1001_g N_A_116_392#_M1004_d VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_369_392#_M1001_d VPB PSHORT L=0.15 W=1
+ AD=0.225 AS=0.175 PD=1.45 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1011 N_A_369_392#_M1011_d N_A2_M1011_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.225 PD=2.59 PS=1.45 NRD=1.9503 NRS=21.67 M=1 R=6.66667
+ SA=75001.8 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__a222oi_1.pxi.spice"
*
.ends
*
*
