* File: sky130_fd_sc_hs__a31oi_1.pxi.spice
* Created: Thu Aug 27 20:29:31 2020
* 
x_PM_SKY130_FD_SC_HS__A31OI_1%A3 N_A3_c_44_n N_A3_M1000_g N_A3_c_45_n
+ N_A3_M1007_g N_A3_c_46_n A3 PM_SKY130_FD_SC_HS__A31OI_1%A3
x_PM_SKY130_FD_SC_HS__A31OI_1%A2 N_A2_c_69_n N_A2_M1005_g N_A2_c_70_n
+ N_A2_M1002_g A2 A2 PM_SKY130_FD_SC_HS__A31OI_1%A2
x_PM_SKY130_FD_SC_HS__A31OI_1%A1 N_A1_c_97_n N_A1_M1001_g N_A1_c_98_n
+ N_A1_M1004_g A1 PM_SKY130_FD_SC_HS__A31OI_1%A1
x_PM_SKY130_FD_SC_HS__A31OI_1%B1 N_B1_M1006_g N_B1_c_133_n N_B1_M1003_g
+ N_B1_c_129_n N_B1_c_130_n B1 B1 N_B1_c_132_n PM_SKY130_FD_SC_HS__A31OI_1%B1
x_PM_SKY130_FD_SC_HS__A31OI_1%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_c_157_n
+ N_VPWR_c_158_n N_VPWR_c_159_n N_VPWR_c_160_n N_VPWR_c_161_n VPWR
+ N_VPWR_c_162_n N_VPWR_c_156_n PM_SKY130_FD_SC_HS__A31OI_1%VPWR
x_PM_SKY130_FD_SC_HS__A31OI_1%A_136_368# N_A_136_368#_M1000_d
+ N_A_136_368#_M1004_d N_A_136_368#_c_193_n N_A_136_368#_c_191_n
+ N_A_136_368#_c_197_n N_A_136_368#_c_201_n N_A_136_368#_c_192_n
+ PM_SKY130_FD_SC_HS__A31OI_1%A_136_368#
x_PM_SKY130_FD_SC_HS__A31OI_1%Y N_Y_M1001_d N_Y_M1003_d N_Y_c_222_n N_Y_c_223_n
+ N_Y_c_224_n N_Y_c_227_n N_Y_c_233_n N_Y_c_225_n Y Y Y N_Y_c_228_n
+ PM_SKY130_FD_SC_HS__A31OI_1%Y
x_PM_SKY130_FD_SC_HS__A31OI_1%VGND N_VGND_M1007_s N_VGND_M1006_d N_VGND_c_278_n
+ N_VGND_c_279_n N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n VGND
+ N_VGND_c_283_n N_VGND_c_284_n PM_SKY130_FD_SC_HS__A31OI_1%VGND
cc_1 VNB N_A3_c_44_n 0.0241262f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.765
cc_2 VNB N_A3_c_45_n 0.0193012f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.22
cc_3 VNB N_A3_c_46_n 0.0564055f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.385
cc_4 VNB A3 0.00839483f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A2_c_69_n 0.0178222f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.765
cc_6 VNB N_A2_c_70_n 0.0376411f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.22
cc_7 VNB A2 0.00485115f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.385
cc_8 VNB N_A1_c_97_n 0.0197655f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.765
cc_9 VNB N_A1_c_98_n 0.0398249f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.22
cc_10 VNB A1 0.00362176f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.385
cc_11 VNB N_B1_c_129_n 0.0206315f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.385
cc_12 VNB N_B1_c_130_n 0.0223503f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_13 VNB B1 0.030738f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_14 VNB N_B1_c_132_n 0.0528453f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_15 VNB N_VPWR_c_156_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_222_n 0.00369921f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.385
cc_17 VNB N_Y_c_223_n 0.00534354f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_Y_c_224_n 6.00478e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_225_n 0.00306185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_278_n 0.0125358f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.385
cc_21 VNB N_VGND_c_279_n 0.0377251f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_VGND_c_280_n 0.0344107f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_23 VNB N_VGND_c_281_n 0.0450666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_282_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_283_n 0.0123263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_284_n 0.19226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_A3_c_44_n 0.0272404f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.765
cc_28 VPB N_A2_c_70_n 0.0234521f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.22
cc_29 VPB N_A1_c_98_n 0.0240609f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.22
cc_30 VPB N_B1_c_133_n 0.0200304f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.22
cc_31 VPB N_B1_c_129_n 0.00895197f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.385
cc_32 VPB N_VPWR_c_157_n 0.0125099f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.385
cc_33 VPB N_VPWR_c_158_n 0.0594617f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_34 VPB N_VPWR_c_159_n 0.00987728f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_35 VPB N_VPWR_c_160_n 0.0212406f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_36 VPB N_VPWR_c_161_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_162_n 0.0384912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_156_n 0.0654951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_136_368#_c_191_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_40 VPB N_A_136_368#_c_192_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_41 VPB N_Y_c_222_n 5.66269e-19 $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.385
cc_42 VPB N_Y_c_227_n 0.0339211f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_43 VPB N_Y_c_228_n 0.0545515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 N_A3_c_45_n N_A2_c_69_n 0.0337327f $X=0.65 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_45 N_A3_c_44_n N_A2_c_70_n 0.0560708f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_46 N_A3_c_45_n A2 8.19586e-19 $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_47 N_A3_c_44_n N_VPWR_c_158_n 0.0337048f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_48 N_A3_c_46_n N_VPWR_c_158_n 0.00245403f $X=0.515 $Y=1.385 $X2=0 $Y2=0
cc_49 A3 N_VPWR_c_158_n 0.0198099f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_A3_c_44_n N_VPWR_c_160_n 0.00445602f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A3_c_44_n N_VPWR_c_156_n 0.00861679f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_52 N_A3_c_44_n N_A_136_368#_c_193_n 0.00208031f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_53 N_A3_c_44_n N_A_136_368#_c_191_n 0.00861647f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_54 N_A3_c_44_n N_Y_c_222_n 0.0180962f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_55 N_A3_c_45_n N_Y_c_222_n 0.0191301f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_56 A3 N_Y_c_222_n 0.0265523f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A3_c_45_n N_Y_c_224_n 0.00539306f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A3_c_44_n N_Y_c_233_n 0.010466f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_59 N_A3_c_45_n N_VGND_c_279_n 0.0179036f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_60 N_A3_c_46_n N_VGND_c_279_n 0.00232901f $X=0.515 $Y=1.385 $X2=0 $Y2=0
cc_61 A3 N_VGND_c_279_n 0.0288422f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A3_c_45_n N_VGND_c_281_n 0.00348163f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A3_c_45_n N_VGND_c_284_n 0.00546242f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_64 N_A2_c_69_n N_A1_c_97_n 0.0265239f $X=1.04 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_65 A2 N_A1_c_97_n 0.00825186f $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_66 N_A2_c_70_n N_A1_c_98_n 0.0492138f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_67 N_A2_c_70_n A1 4.06701e-19 $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_68 A2 A1 0.0242365f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_69 N_A2_c_70_n N_VPWR_c_159_n 0.00909103f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A2_c_70_n N_VPWR_c_160_n 0.00445602f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A2_c_70_n N_VPWR_c_156_n 0.00859428f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A2_c_70_n N_A_136_368#_c_193_n 4.27055e-19 $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A2_c_70_n N_A_136_368#_c_191_n 0.010066f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A2_c_70_n N_A_136_368#_c_197_n 0.0127987f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A2_c_70_n N_A_136_368#_c_192_n 8.55427e-19 $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A2_c_69_n N_Y_c_222_n 0.0133177f $X=1.04 $Y=1.22 $X2=0 $Y2=0
cc_77 A2 N_Y_c_222_n 0.0554335f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_78 N_A2_c_69_n N_Y_c_223_n 0.0109398f $X=1.04 $Y=1.22 $X2=0 $Y2=0
cc_79 A2 N_Y_c_223_n 0.013653f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A2_c_70_n N_Y_c_227_n 0.0134331f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_81 A2 N_Y_c_227_n 0.0272275f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_82 N_A2_c_69_n N_VGND_c_281_n 0.00291649f $X=1.04 $Y=1.22 $X2=0 $Y2=0
cc_83 N_A2_c_69_n N_VGND_c_284_n 0.00359136f $X=1.04 $Y=1.22 $X2=0 $Y2=0
cc_84 A2 A_223_74# 0.00606047f $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_85 N_A1_c_98_n N_B1_c_133_n 0.0246103f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A1_c_98_n N_B1_c_129_n 0.0270818f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_87 A1 N_B1_c_129_n 3.68035e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A1_c_97_n N_B1_c_130_n 0.0233894f $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_89 N_A1_c_98_n B1 0.00216087f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_90 A1 B1 0.029889f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A1_c_98_n N_VPWR_c_159_n 0.00902378f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A1_c_98_n N_VPWR_c_162_n 0.00445602f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A1_c_98_n N_VPWR_c_156_n 0.00860083f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A1_c_98_n N_A_136_368#_c_191_n 8.50228e-19 $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A1_c_98_n N_A_136_368#_c_197_n 0.0127987f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A1_c_98_n N_A_136_368#_c_201_n 4.27055e-19 $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A1_c_98_n N_A_136_368#_c_192_n 0.0102039f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A1_c_97_n N_Y_c_223_n 0.0131896f $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_99 A1 N_Y_c_223_n 0.00420927f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A1_c_98_n N_Y_c_227_n 0.013694f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_101 A1 N_Y_c_227_n 0.024317f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_102 N_A1_c_98_n N_Y_c_225_n 9.02817e-19 $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_103 A1 N_Y_c_225_n 0.0111615f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A1_c_98_n N_Y_c_228_n 7.47851e-19 $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A1_c_97_n N_VGND_c_280_n 7.24629e-19 $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A1_c_97_n N_VGND_c_281_n 0.00291649f $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A1_c_97_n N_VGND_c_284_n 0.00361625f $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_108 N_B1_c_133_n N_VPWR_c_162_n 0.00445602f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_109 N_B1_c_133_n N_VPWR_c_156_n 0.00862822f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_110 N_B1_c_133_n N_A_136_368#_c_192_n 0.00405513f $X=2.195 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_B1_c_133_n N_Y_c_227_n 0.010996f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_112 N_B1_c_129_n N_Y_c_227_n 0.00541994f $X=2.285 $Y=1.385 $X2=0 $Y2=0
cc_113 B1 N_Y_c_227_n 0.0579042f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B1_c_132_n N_Y_c_227_n 0.0109287f $X=2.61 $Y=1.385 $X2=0 $Y2=0
cc_115 N_B1_c_130_n N_Y_c_225_n 0.00110948f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_116 B1 N_Y_c_225_n 7.29591e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B1_c_133_n N_Y_c_228_n 0.0137364f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_118 N_B1_c_129_n N_VGND_c_280_n 0.00199643f $X=2.285 $Y=1.385 $X2=0 $Y2=0
cc_119 N_B1_c_130_n N_VGND_c_280_n 0.0124734f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_120 B1 N_VGND_c_280_n 0.0259403f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_121 N_B1_c_130_n N_VGND_c_281_n 0.00383152f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_122 N_B1_c_130_n N_VGND_c_284_n 0.00758792f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_123 N_VPWR_c_158_n N_A_136_368#_c_193_n 0.0118923f $X=0.29 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_VPWR_c_158_n N_A_136_368#_c_191_n 0.0494855f $X=0.29 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_VPWR_c_159_n N_A_136_368#_c_191_n 0.0383004f $X=1.37 $Y=2.485 $X2=0
+ $Y2=0
cc_126 N_VPWR_c_160_n N_A_136_368#_c_191_n 0.014552f $X=1.205 $Y=3.33 $X2=0
+ $Y2=0
cc_127 N_VPWR_c_156_n N_A_136_368#_c_191_n 0.0119791f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_128 N_VPWR_M1002_d N_A_136_368#_c_197_n 0.0103777f $X=1.13 $Y=1.84 $X2=0
+ $Y2=0
cc_129 N_VPWR_c_159_n N_A_136_368#_c_197_n 0.0266856f $X=1.37 $Y=2.485 $X2=0
+ $Y2=0
cc_130 N_VPWR_c_159_n N_A_136_368#_c_192_n 0.0369621f $X=1.37 $Y=2.485 $X2=0
+ $Y2=0
cc_131 N_VPWR_c_162_n N_A_136_368#_c_192_n 0.0145938f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_132 N_VPWR_c_156_n N_A_136_368#_c_192_n 0.0120466f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_133 N_VPWR_M1002_d N_Y_c_227_n 0.00427791f $X=1.13 $Y=1.84 $X2=0 $Y2=0
cc_134 N_VPWR_c_158_n N_Y_c_233_n 0.00579827f $X=0.29 $Y=1.985 $X2=0 $Y2=0
cc_135 N_VPWR_c_162_n N_Y_c_228_n 0.0221794f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_136 N_VPWR_c_156_n N_Y_c_228_n 0.0183253f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_137 N_A_136_368#_M1000_d N_Y_c_227_n 0.00135003f $X=0.68 $Y=1.84 $X2=0 $Y2=0
cc_138 N_A_136_368#_M1004_d N_Y_c_227_n 0.00250873f $X=1.77 $Y=1.84 $X2=0 $Y2=0
cc_139 N_A_136_368#_c_193_n N_Y_c_227_n 0.0114779f $X=0.83 $Y=2.23 $X2=0 $Y2=0
cc_140 N_A_136_368#_c_197_n N_Y_c_227_n 0.045543f $X=1.755 $Y=2.145 $X2=0 $Y2=0
cc_141 N_A_136_368#_c_201_n N_Y_c_227_n 0.0203011f $X=1.92 $Y=2.23 $X2=0 $Y2=0
cc_142 N_A_136_368#_M1000_d N_Y_c_233_n 6.41842e-19 $X=0.68 $Y=1.84 $X2=0 $Y2=0
cc_143 N_A_136_368#_c_193_n N_Y_c_233_n 0.00645682f $X=0.83 $Y=2.23 $X2=0 $Y2=0
cc_144 N_A_136_368#_c_192_n N_Y_c_228_n 0.0307786f $X=1.92 $Y=2.825 $X2=0 $Y2=0
cc_145 N_Y_c_222_n N_VGND_c_279_n 0.0362227f $X=0.71 $Y=1.72 $X2=0 $Y2=0
cc_146 N_Y_c_224_n N_VGND_c_279_n 0.0140387f $X=0.795 $Y=0.435 $X2=0 $Y2=0
cc_147 N_Y_c_225_n N_VGND_c_280_n 0.00729487f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_148 N_Y_c_223_n N_VGND_c_281_n 0.0369511f $X=1.73 $Y=0.435 $X2=0 $Y2=0
cc_149 N_Y_c_224_n N_VGND_c_281_n 0.00728664f $X=0.795 $Y=0.435 $X2=0 $Y2=0
cc_150 N_Y_c_225_n N_VGND_c_281_n 0.014693f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_151 N_Y_c_223_n N_VGND_c_284_n 0.0316226f $X=1.73 $Y=0.435 $X2=0 $Y2=0
cc_152 N_Y_c_224_n N_VGND_c_284_n 0.00579633f $X=0.795 $Y=0.435 $X2=0 $Y2=0
cc_153 N_Y_c_225_n N_VGND_c_284_n 0.0121757f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_154 N_Y_c_222_n A_145_74# 0.00586266f $X=0.71 $Y=1.72 $X2=-0.19 $Y2=-0.245
cc_155 N_Y_c_223_n A_145_74# 0.00427342f $X=1.73 $Y=0.435 $X2=-0.19 $Y2=-0.245
cc_156 N_Y_c_223_n A_223_74# 0.00868086f $X=1.73 $Y=0.435 $X2=-0.19 $Y2=-0.245
