* File: sky130_fd_sc_hs__o221a_2.spice
* Created: Tue Sep  1 20:15:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o221a_2.pex.spice"
.subckt sky130_fd_sc_hs__o221a_2  VNB VPB C1 B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1006 N_A_165_74#_M1006_d N_C1_M1006_g N_A_27_368#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.12765 AS=0.2109 PD=1.085 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_264_74#_M1010_d N_B1_M1010_g N_A_165_74#_M1006_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.13135 AS=0.12765 PD=1.095 PS=1.085 NRD=5.664 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_A_165_74#_M1003_d N_B2_M1003_g N_A_264_74#_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.13135 PD=2.05 PS=1.095 NRD=0 NRS=6.48 M=1 R=4.93333
+ SA=75001.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_264_74#_M1012_d N_A2_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_264_74#_M1012_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1004_d N_A_27_368#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_27_368#_M1007_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3108 AS=0.1036 PD=2.32 PS=1.02 NRD=21.888 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1013 N_VPWR_M1013_d N_C1_M1013_g N_A_27_368#_M1013_s VPB PSHORT L=0.15 W=1
+ AD=0.465 AS=0.295 PD=1.93 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75004 A=0.15 P=2.3 MULT=1
MM1002 A_332_368# N_B1_M1002_g N_VPWR_M1013_d VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.465 PD=1.27 PS=1.93 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75001.3
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1008 N_A_27_368#_M1008_d N_B2_M1008_g A_332_368# VPB PSHORT L=0.15 W=1 AD=0.21
+ AS=0.135 PD=1.42 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75001.7
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1011 A_530_368# N_A2_M1011_g N_A_27_368#_M1008_d VPB PSHORT L=0.15 W=1 AD=0.21
+ AS=0.21 PD=1.42 PS=1.42 NRD=30.5153 NRS=25.5903 M=1 R=6.66667 SA=75002.3
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_530_368# VPB PSHORT L=0.15 W=1 AD=0.278962
+ AS=0.21 PD=1.57547 PS=1.42 NRD=41.8428 NRS=30.5153 M=1 R=6.66667 SA=75002.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_27_368#_M1001_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.312438 PD=1.42 PS=1.76453 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1005 N_X_M1001_d N_A_27_368#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_hs__o221a_2.pxi.spice"
*
.ends
*
*
