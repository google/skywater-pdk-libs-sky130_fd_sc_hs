# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__o21bai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21bai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 3.715000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.450000 7.075000 1.780000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.855000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.370000 1.950000 5.625000 2.020000 ;
        RECT 2.370000 2.020000 4.710000 2.120000 ;
        RECT 2.370000 2.120000 2.620000 2.735000 ;
        RECT 3.320000 2.120000 3.650000 2.735000 ;
        RECT 3.965000 1.010000 5.595000 1.180000 ;
        RECT 3.965000 1.180000 4.195000 1.950000 ;
        RECT 4.265000 0.595000 4.595000 1.010000 ;
        RECT 4.380000 1.850000 5.625000 1.950000 ;
        RECT 4.380000 2.120000 4.710000 2.980000 ;
        RECT 5.265000 0.595000 5.595000 1.010000 ;
        RECT 5.295000 2.020000 5.625000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 3.075000 1.180000 ;
      RECT 0.120000  1.950000 2.170000 2.120000 ;
      RECT 0.120000  2.120000 0.370000 2.980000 ;
      RECT 0.545000  0.085000 0.875000 0.840000 ;
      RECT 0.570000  2.290000 0.820000 3.245000 ;
      RECT 1.020000  2.120000 1.270000 2.980000 ;
      RECT 1.105000  0.350000 1.275000 1.010000 ;
      RECT 1.455000  0.085000 1.785000 0.840000 ;
      RECT 1.470000  2.290000 1.800000 3.245000 ;
      RECT 1.965000  0.350000 2.135000 1.010000 ;
      RECT 2.000000  1.820000 2.170000 1.950000 ;
      RECT 2.000000  2.120000 2.170000 2.905000 ;
      RECT 2.000000  2.905000 4.150000 3.075000 ;
      RECT 2.315000  0.085000 2.645000 0.840000 ;
      RECT 2.820000  2.290000 3.150000 2.905000 ;
      RECT 2.825000  0.350000 3.075000 0.670000 ;
      RECT 2.825000  0.670000 4.095000 0.840000 ;
      RECT 2.825000  0.840000 3.075000 1.010000 ;
      RECT 3.255000  0.085000 3.585000 0.500000 ;
      RECT 3.765000  0.255000 6.095000 0.425000 ;
      RECT 3.765000  0.425000 4.095000 0.670000 ;
      RECT 3.820000  2.290000 4.150000 2.905000 ;
      RECT 4.370000  1.350000 5.965000 1.680000 ;
      RECT 4.765000  0.425000 5.095000 0.840000 ;
      RECT 4.910000  2.190000 5.080000 3.245000 ;
      RECT 5.765000  0.425000 6.095000 0.940000 ;
      RECT 5.795000  1.110000 6.575000 1.280000 ;
      RECT 5.795000  1.280000 5.965000 1.350000 ;
      RECT 5.795000  1.680000 5.965000 1.950000 ;
      RECT 5.795000  1.950000 6.555000 2.120000 ;
      RECT 5.855000  2.290000 6.105000 3.245000 ;
      RECT 6.305000  2.120000 6.555000 2.980000 ;
      RECT 6.325000  0.500000 6.575000 1.110000 ;
      RECT 6.755000  0.085000 7.085000 1.280000 ;
      RECT 6.755000  2.100000 7.085000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__o21bai_4
END LIBRARY
