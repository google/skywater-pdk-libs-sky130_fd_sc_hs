* File: sky130_fd_sc_hs__nand2b_4.spice
* Created: Tue Sep  1 20:09:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nand2b_4.pex.spice"
.subckt sky130_fd_sc_hs__nand2b_4  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_N_M1012_g N_A_31_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_31_74#_M1000_g N_A_243_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.9 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1000_d N_A_31_74#_M1007_g N_A_243_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1010_d N_A_31_74#_M1010_g N_A_243_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.15355 AS=0.1036 PD=1.155 PS=1.02 NRD=12.156 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75003 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1010_d N_A_31_74#_M1014_g N_A_243_74#_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.15355 AS=0.1036 PD=1.155 PS=1.02 NRD=9.72 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1001 N_A_243_74#_M1014_s N_B_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1004 N_A_243_74#_M1004_d N_B_M1004_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1009 N_A_243_74#_M1004_d N_B_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.27935 PD=1.02 PS=1.495 NRD=0 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_A_243_74#_M1011_d N_B_M1011_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.27935 PD=2.05 PS=1.495 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_31_74#_M1005_d N_A_N_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.5376 PD=1.14 PS=2.96 NRD=2.3443 NRS=3.5066 M=1 R=5.6 SA=75000.6
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1008 N_A_31_74#_M1005_d N_A_N_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.174 PD=1.14 PS=1.29 NRD=2.3443 NRS=22.261 M=1 R=5.6 SA=75001
+ SB=75003.8 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_31_74#_M1003_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3808 AS=0.232 PD=1.8 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75003.3 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1003_d N_A_31_74#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3808 AS=0.896 PD=1.8 PS=2.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75002.4 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1006_s N_B_M1002_g N_Y_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.896
+ AS=0.1792 PD=2.72 PS=1.44 NRD=7.0329 NRS=5.2599 M=1 R=7.46667 SA=75003.8
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_B_M1013_g N_Y_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.336
+ AS=0.1792 PD=2.84 PS=1.44 NRD=2.6201 NRS=1.7533 M=1 R=7.46667 SA=75004.3
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX15_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_hs__nand2b_4.pxi.spice"
*
.ends
*
*
