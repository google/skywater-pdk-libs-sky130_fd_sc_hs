* File: sky130_fd_sc_hs__a32oi_4.pex.spice
* Created: Thu Aug 27 20:30:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A32OI_4%B2 3 5 7 10 12 14 17 19 21 22 24 27 29 30 31
+ 32 49
c79 27 0 8.12065e-20 $X=1.92 $Y=0.74
c80 22 0 1.39988e-19 $X=1.905 $Y=1.765
r81 49 50 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=1.905 $Y=1.557
+ $X2=1.92 $Y2=1.557
r82 47 49 39.2935 $w=3.68e-07 $l=3e-07 $layer=POLY_cond $X=1.605 $Y=1.557
+ $X2=1.905 $Y2=1.557
r83 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.605
+ $Y=1.515 $X2=1.605 $Y2=1.515
r84 45 47 19.6467 $w=3.68e-07 $l=1.5e-07 $layer=POLY_cond $X=1.455 $Y=1.557
+ $X2=1.605 $Y2=1.557
r85 44 45 3.92935 $w=3.68e-07 $l=3e-08 $layer=POLY_cond $X=1.425 $Y=1.557
+ $X2=1.455 $Y2=1.557
r86 43 44 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=1.005 $Y=1.557
+ $X2=1.425 $Y2=1.557
r87 42 43 1.30978 $w=3.68e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.557
+ $X2=1.005 $Y2=1.557
r88 40 42 53.7011 $w=3.68e-07 $l=4.1e-07 $layer=POLY_cond $X=0.585 $Y=1.557
+ $X2=0.995 $Y2=1.557
r89 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r90 38 40 9.82337 $w=3.68e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.585 $Y2=1.557
r91 37 38 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r92 32 48 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.605 $Y2=1.565
r93 31 48 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.605 $Y2=1.565
r94 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r95 30 41 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r96 29 41 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r97 25 50 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.92 $Y=1.35
+ $X2=1.92 $Y2=1.557
r98 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.92 $Y=1.35
+ $X2=1.92 $Y2=0.74
r99 22 49 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=1.557
r100 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=2.4
r101 19 45 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.557
r102 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r103 15 44 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.557
r104 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.74
r105 12 43 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.557
r106 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r107 8 42 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.557
r108 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r109 5 38 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r110 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r111 1 37 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r112 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%B1 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 33 50
c90 33 0 2.03596e-19 $X=4.08 $Y=1.665
c91 26 0 4.35069e-20 $X=3.905 $Y=1.765
c92 17 0 8.60869e-20 $X=3.28 $Y=0.74
c93 3 0 7.59056e-20 $X=2.35 $Y=0.74
r94 50 52 13.8658 $w=3.65e-07 $l=1.05e-07 $layer=POLY_cond $X=3.8 $Y=1.557
+ $X2=3.905 $Y2=1.557
r95 50 51 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.8
+ $Y=1.515 $X2=3.8 $Y2=1.515
r96 48 50 11.8849 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=3.71 $Y=1.557 $X2=3.8
+ $Y2=1.557
r97 47 48 40.2767 $w=3.65e-07 $l=3.05e-07 $layer=POLY_cond $X=3.405 $Y=1.557
+ $X2=3.71 $Y2=1.557
r98 46 47 16.5068 $w=3.65e-07 $l=1.25e-07 $layer=POLY_cond $X=3.28 $Y=1.557
+ $X2=3.405 $Y2=1.557
r99 45 46 49.5205 $w=3.65e-07 $l=3.75e-07 $layer=POLY_cond $X=2.905 $Y=1.557
+ $X2=3.28 $Y2=1.557
r100 44 45 16.5068 $w=3.65e-07 $l=1.25e-07 $layer=POLY_cond $X=2.78 $Y=1.557
+ $X2=2.905 $Y2=1.557
r101 42 44 44.8986 $w=3.65e-07 $l=3.4e-07 $layer=POLY_cond $X=2.44 $Y=1.557
+ $X2=2.78 $Y2=1.557
r102 42 43 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.44
+ $Y=1.515 $X2=2.44 $Y2=1.515
r103 40 42 4.62192 $w=3.65e-07 $l=3.5e-08 $layer=POLY_cond $X=2.405 $Y=1.557
+ $X2=2.44 $Y2=1.557
r104 39 40 7.26301 $w=3.65e-07 $l=5.5e-08 $layer=POLY_cond $X=2.35 $Y=1.557
+ $X2=2.405 $Y2=1.557
r105 33 51 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.8 $Y2=1.565
r106 32 51 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.8
+ $Y2=1.565
r107 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r108 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r109 30 43 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.44
+ $Y2=1.565
r110 29 43 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.44 $Y2=1.565
r111 26 52 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.905 $Y=1.765
+ $X2=3.905 $Y2=1.557
r112 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.905 $Y=1.765
+ $X2=3.905 $Y2=2.4
r113 22 48 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=1.557
r114 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=0.74
r115 19 47 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=1.557
r116 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=2.4
r117 15 46 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.28 $Y=1.35
+ $X2=3.28 $Y2=1.557
r118 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.28 $Y=1.35
+ $X2=3.28 $Y2=0.74
r119 12 45 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.905 $Y=1.765
+ $X2=2.905 $Y2=1.557
r120 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.905 $Y=1.765
+ $X2=2.905 $Y2=2.4
r121 8 44 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.78 $Y=1.35
+ $X2=2.78 $Y2=1.557
r122 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.78 $Y=1.35
+ $X2=2.78 $Y2=0.74
r123 5 40 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.557
r124 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r125 1 39 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=1.35
+ $X2=2.35 $Y2=1.557
r126 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.35 $Y=1.35 $X2=2.35
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 46 47
c81 46 0 4.35069e-20 $X=5.64 $Y=1.515
c82 1 0 6.36075e-20 $X=4.545 $Y=1.765
r83 47 48 1.97541 $w=3.66e-07 $l=1.5e-08 $layer=POLY_cond $X=6.045 $Y=1.557
+ $X2=6.06 $Y2=1.557
r84 45 47 53.3361 $w=3.66e-07 $l=4.05e-07 $layer=POLY_cond $X=5.64 $Y=1.557
+ $X2=6.045 $Y2=1.557
r85 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.64
+ $Y=1.515 $X2=5.64 $Y2=1.515
r86 43 45 1.31694 $w=3.66e-07 $l=1e-08 $layer=POLY_cond $X=5.63 $Y=1.557
+ $X2=5.64 $Y2=1.557
r87 42 43 17.7787 $w=3.66e-07 $l=1.35e-07 $layer=POLY_cond $X=5.495 $Y=1.557
+ $X2=5.63 $Y2=1.557
r88 41 42 38.8497 $w=3.66e-07 $l=2.95e-07 $layer=POLY_cond $X=5.2 $Y=1.557
+ $X2=5.495 $Y2=1.557
r89 40 41 20.4126 $w=3.66e-07 $l=1.55e-07 $layer=POLY_cond $X=5.045 $Y=1.557
+ $X2=5.2 $Y2=1.557
r90 39 40 45.4344 $w=3.66e-07 $l=3.45e-07 $layer=POLY_cond $X=4.7 $Y=1.557
+ $X2=5.045 $Y2=1.557
r91 37 39 10.5355 $w=3.66e-07 $l=8e-08 $layer=POLY_cond $X=4.62 $Y=1.557 $X2=4.7
+ $Y2=1.557
r92 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.62
+ $Y=1.515 $X2=4.62 $Y2=1.515
r93 35 37 9.87705 $w=3.66e-07 $l=7.5e-08 $layer=POLY_cond $X=4.545 $Y=1.557
+ $X2=4.62 $Y2=1.557
r94 31 46 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.64 $Y2=1.565
r95 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r96 30 38 11.2564 $w=4.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.62 $Y2=1.565
r97 29 38 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=4.56 $Y=1.565 $X2=4.62
+ $Y2=1.565
r98 25 48 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.06 $Y=1.35
+ $X2=6.06 $Y2=1.557
r99 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.06 $Y=1.35
+ $X2=6.06 $Y2=0.74
r100 22 47 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.045 $Y=1.765
+ $X2=6.045 $Y2=1.557
r101 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.045 $Y=1.765
+ $X2=6.045 $Y2=2.4
r102 18 43 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.63 $Y=1.35
+ $X2=5.63 $Y2=1.557
r103 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.63 $Y=1.35
+ $X2=5.63 $Y2=0.74
r104 15 42 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.495 $Y=1.765
+ $X2=5.495 $Y2=1.557
r105 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.495 $Y=1.765
+ $X2=5.495 $Y2=2.4
r106 11 41 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.2 $Y=1.35
+ $X2=5.2 $Y2=1.557
r107 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.2 $Y=1.35 $X2=5.2
+ $Y2=0.74
r108 8 40 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.045 $Y=1.765
+ $X2=5.045 $Y2=1.557
r109 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.045 $Y=1.765
+ $X2=5.045 $Y2=2.4
r110 4 39 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.7 $Y=1.35 $X2=4.7
+ $Y2=1.557
r111 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.7 $Y=1.35 $X2=4.7
+ $Y2=0.74
r112 1 35 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.545 $Y=1.765
+ $X2=4.545 $Y2=1.557
r113 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.545 $Y=1.765
+ $X2=4.545 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%A2 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 48
c90 48 0 1.89024e-19 $X=7.92 $Y=1.515
c91 32 0 1.23692e-20 $X=8.4 $Y=1.665
c92 26 0 1.28414e-19 $X=7.995 $Y=1.765
c93 5 0 6.40318e-20 $X=6.505 $Y=1.765
r94 48 50 9.87705 $w=3.66e-07 $l=7.5e-08 $layer=POLY_cond $X=7.92 $Y=1.557
+ $X2=7.995 $Y2=1.557
r95 46 48 17.7787 $w=3.66e-07 $l=1.35e-07 $layer=POLY_cond $X=7.785 $Y=1.557
+ $X2=7.92 $Y2=1.557
r96 45 46 38.1913 $w=3.66e-07 $l=2.9e-07 $layer=POLY_cond $X=7.495 $Y=1.557
+ $X2=7.785 $Y2=1.557
r97 44 45 18.4372 $w=3.66e-07 $l=1.4e-07 $layer=POLY_cond $X=7.355 $Y=1.557
+ $X2=7.495 $Y2=1.557
r98 43 44 40.8251 $w=3.66e-07 $l=3.1e-07 $layer=POLY_cond $X=7.045 $Y=1.557
+ $X2=7.355 $Y2=1.557
r99 42 43 16.4617 $w=3.66e-07 $l=1.25e-07 $layer=POLY_cond $X=6.92 $Y=1.557
+ $X2=7.045 $Y2=1.557
r100 40 42 2.63388 $w=3.66e-07 $l=2e-08 $layer=POLY_cond $X=6.9 $Y=1.557
+ $X2=6.92 $Y2=1.557
r101 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.9
+ $Y=1.515 $X2=6.9 $Y2=1.515
r102 38 40 52.0191 $w=3.66e-07 $l=3.95e-07 $layer=POLY_cond $X=6.505 $Y=1.557
+ $X2=6.9 $Y2=1.557
r103 37 38 1.97541 $w=3.66e-07 $l=1.5e-08 $layer=POLY_cond $X=6.49 $Y=1.557
+ $X2=6.505 $Y2=1.557
r104 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.4 $Y2=1.565
r105 31 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.92
+ $Y=1.515 $X2=7.92 $Y2=1.515
r106 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r107 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r108 29 41 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=6.96 $Y=1.565 $X2=6.9
+ $Y2=1.565
r109 26 50 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.995 $Y=1.765
+ $X2=7.995 $Y2=1.557
r110 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.995 $Y=1.765
+ $X2=7.995 $Y2=2.4
r111 22 46 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.785 $Y=1.35
+ $X2=7.785 $Y2=1.557
r112 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.785 $Y=1.35
+ $X2=7.785 $Y2=0.74
r113 19 45 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.495 $Y=1.765
+ $X2=7.495 $Y2=1.557
r114 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.495 $Y=1.765
+ $X2=7.495 $Y2=2.4
r115 15 44 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.355 $Y=1.35
+ $X2=7.355 $Y2=1.557
r116 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.355 $Y=1.35
+ $X2=7.355 $Y2=0.74
r117 12 43 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.045 $Y=1.765
+ $X2=7.045 $Y2=1.557
r118 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.045 $Y=1.765
+ $X2=7.045 $Y2=2.4
r119 8 42 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.92 $Y=1.35
+ $X2=6.92 $Y2=1.557
r120 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.92 $Y=1.35
+ $X2=6.92 $Y2=0.74
r121 5 38 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.505 $Y=1.765
+ $X2=6.505 $Y2=1.557
r122 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.505 $Y=1.765
+ $X2=6.505 $Y2=2.4
r123 1 37 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.49 $Y=1.35
+ $X2=6.49 $Y2=1.557
r124 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.49 $Y=1.35 $X2=6.49
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 49
c84 32 0 1.89024e-19 $X=10.32 $Y=1.665
c85 8 0 1.23692e-20 $X=8.995 $Y=1.765
r86 49 50 2.16467 $w=3.34e-07 $l=1.5e-08 $layer=POLY_cond $X=10.05 $Y=1.557
+ $X2=10.065 $Y2=1.557
r87 47 49 14.4311 $w=3.34e-07 $l=1e-07 $layer=POLY_cond $X=9.95 $Y=1.557
+ $X2=10.05 $Y2=1.557
r88 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.95
+ $Y=1.515 $X2=9.95 $Y2=1.515
r89 45 47 45.4581 $w=3.34e-07 $l=3.15e-07 $layer=POLY_cond $X=9.635 $Y=1.557
+ $X2=9.95 $Y2=1.557
r90 44 45 20.2036 $w=3.34e-07 $l=1.4e-07 $layer=POLY_cond $X=9.495 $Y=1.557
+ $X2=9.635 $Y2=1.557
r91 42 44 32.4701 $w=3.34e-07 $l=2.25e-07 $layer=POLY_cond $X=9.27 $Y=1.557
+ $X2=9.495 $Y2=1.557
r92 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.27
+ $Y=1.515 $X2=9.27 $Y2=1.515
r93 40 42 9.38024 $w=3.34e-07 $l=6.5e-08 $layer=POLY_cond $X=9.205 $Y=1.557
+ $X2=9.27 $Y2=1.557
r94 39 40 30.3054 $w=3.34e-07 $l=2.1e-07 $layer=POLY_cond $X=8.995 $Y=1.557
+ $X2=9.205 $Y2=1.557
r95 38 39 31.7485 $w=3.34e-07 $l=2.2e-07 $layer=POLY_cond $X=8.775 $Y=1.557
+ $X2=8.995 $Y2=1.557
r96 37 38 40.4072 $w=3.34e-07 $l=2.8e-07 $layer=POLY_cond $X=8.495 $Y=1.557
+ $X2=8.775 $Y2=1.557
r97 32 48 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=9.95 $Y2=1.565
r98 31 48 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.95 $Y2=1.565
r99 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.84 $Y2=1.565
r100 30 43 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.27 $Y2=1.565
r101 29 43 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.27 $Y2=1.565
r102 25 50 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.065 $Y=1.35
+ $X2=10.065 $Y2=1.557
r103 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.065 $Y=1.35
+ $X2=10.065 $Y2=0.74
r104 22 49 21.5099 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.05 $Y=1.765
+ $X2=10.05 $Y2=1.557
r105 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.05 $Y=1.765
+ $X2=10.05 $Y2=2.4
r106 18 45 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.635 $Y=1.35
+ $X2=9.635 $Y2=1.557
r107 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.635 $Y=1.35
+ $X2=9.635 $Y2=0.74
r108 15 44 21.5099 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.495 $Y=1.765
+ $X2=9.495 $Y2=1.557
r109 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.495 $Y=1.765
+ $X2=9.495 $Y2=2.4
r110 11 40 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.205 $Y=1.35
+ $X2=9.205 $Y2=1.557
r111 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.205 $Y=1.35
+ $X2=9.205 $Y2=0.74
r112 8 39 21.5099 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.995 $Y=1.765
+ $X2=8.995 $Y2=1.557
r113 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.995 $Y=1.765
+ $X2=8.995 $Y2=2.4
r114 4 38 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.775 $Y=1.35
+ $X2=8.775 $Y2=1.557
r115 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.775 $Y=1.35
+ $X2=8.775 $Y2=0.74
r116 1 37 21.5099 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.495 $Y=1.765
+ $X2=8.495 $Y2=1.557
r117 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.495 $Y=1.765
+ $X2=8.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%A_27_368# 1 2 3 4 5 6 7 8 9 10 11 36 40 41
+ 44 46 50 52 56 58 60 61 62 66 70 72 73 76 78 82 84 88 90 92 94 96 97 98 102
+ 104 107 109 111
c172 104 0 6.40318e-20 $X=6.27 $Y=2.455
c173 76 0 1.28414e-19 $X=7.27 $Y=2.815
r174 92 113 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=2.12
+ $X2=10.275 $Y2=2.035
r175 92 94 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=10.275 $Y=2.12
+ $X2=10.275 $Y2=2.815
r176 91 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=2.035
+ $X2=9.27 $Y2=2.035
r177 90 113 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.11 $Y=2.035
+ $X2=10.275 $Y2=2.035
r178 90 91 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=10.11 $Y=2.035
+ $X2=9.435 $Y2=2.035
r179 86 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.27 $Y=2.12
+ $X2=9.27 $Y2=2.035
r180 86 88 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.27 $Y=2.12
+ $X2=9.27 $Y2=2.815
r181 85 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.435 $Y=2.035
+ $X2=8.27 $Y2=2.035
r182 84 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=2.035
+ $X2=9.27 $Y2=2.035
r183 84 85 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.105 $Y=2.035
+ $X2=8.435 $Y2=2.035
r184 80 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.27 $Y=2.12
+ $X2=8.27 $Y2=2.035
r185 80 82 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.27 $Y=2.12
+ $X2=8.27 $Y2=2.815
r186 79 106 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=2.035
+ $X2=7.27 $Y2=2.035
r187 78 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.105 $Y=2.035
+ $X2=8.27 $Y2=2.035
r188 78 79 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.105 $Y=2.035
+ $X2=7.435 $Y2=2.035
r189 74 107 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.27 $Y=2.46
+ $X2=7.27 $Y2=2.375
r190 74 76 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.27 $Y=2.46
+ $X2=7.27 $Y2=2.815
r191 73 107 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.27 $Y=2.29
+ $X2=7.27 $Y2=2.375
r192 72 106 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.27 $Y=2.12
+ $X2=7.27 $Y2=2.035
r193 72 73 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.27 $Y=2.12
+ $X2=7.27 $Y2=2.29
r194 71 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=2.375
+ $X2=6.27 $Y2=2.375
r195 70 107 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.105 $Y=2.375
+ $X2=7.27 $Y2=2.375
r196 70 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.105 $Y=2.375
+ $X2=6.435 $Y2=2.375
r197 67 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=2.375
+ $X2=5.27 $Y2=2.375
r198 66 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=2.375
+ $X2=6.27 $Y2=2.375
r199 66 67 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.105 $Y=2.375
+ $X2=5.435 $Y2=2.375
r200 63 100 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=2.375
+ $X2=4.18 $Y2=2.375
r201 62 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.105 $Y=2.375
+ $X2=5.27 $Y2=2.375
r202 62 63 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.105 $Y=2.375
+ $X2=4.345 $Y2=2.375
r203 60 100 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=2.46
+ $X2=4.18 $Y2=2.375
r204 60 61 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.18 $Y=2.46
+ $X2=4.18 $Y2=2.905
r205 59 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=2.99
+ $X2=3.18 $Y2=2.99
r206 58 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.015 $Y=2.99
+ $X2=4.18 $Y2=2.905
r207 58 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.015 $Y=2.99
+ $X2=3.345 $Y2=2.99
r208 54 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=2.905
+ $X2=3.18 $Y2=2.99
r209 54 56 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.18 $Y=2.905
+ $X2=3.18 $Y2=2.455
r210 53 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=2.99
+ $X2=2.18 $Y2=2.99
r211 52 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=2.99
+ $X2=3.18 $Y2=2.99
r212 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.015 $Y=2.99
+ $X2=2.345 $Y2=2.99
r213 48 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.905
+ $X2=2.18 $Y2=2.99
r214 48 50 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.18 $Y=2.905
+ $X2=2.18 $Y2=2.455
r215 47 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.99
+ $X2=1.23 $Y2=2.99
r216 46 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=2.18 $Y2=2.99
r217 46 47 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=1.315 $Y2=2.99
r218 42 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.99
r219 42 44 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.455
r220 40 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=1.23 $Y2=2.99
r221 40 41 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=0.445 $Y2=2.99
r222 36 39 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r223 34 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r224 34 39 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r225 11 113 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=10.125
+ $Y=1.84 $X2=10.275 $Y2=2.115
r226 11 94 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.125
+ $Y=1.84 $X2=10.275 $Y2=2.815
r227 10 111 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=9.07
+ $Y=1.84 $X2=9.27 $Y2=2.115
r228 10 88 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=9.07
+ $Y=1.84 $X2=9.27 $Y2=2.815
r229 9 109 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=1.84 $X2=8.27 $Y2=2.115
r230 9 82 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=1.84 $X2=8.27 $Y2=2.815
r231 8 106 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=7.12
+ $Y=1.84 $X2=7.27 $Y2=2.115
r232 8 76 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.12
+ $Y=1.84 $X2=7.27 $Y2=2.815
r233 7 104 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.12
+ $Y=1.84 $X2=6.27 $Y2=2.455
r234 6 102 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.12
+ $Y=1.84 $X2=5.27 $Y2=2.455
r235 5 100 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=3.98
+ $Y=1.84 $X2=4.18 $Y2=2.455
r236 4 56 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=2.98
+ $Y=1.84 $X2=3.18 $Y2=2.455
r237 3 50 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=1.98
+ $Y=1.84 $X2=2.18 $Y2=2.455
r238 2 44 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=2.455
r239 1 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r240 1 36 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%Y 1 2 3 4 5 6 7 8 27 31 35 39 45 48 50 52 54
+ 59 60 62 63 64 65 66 79 81
c125 54 0 8.12065e-20 $X=2.565 $Y=0.86
c126 35 0 7.59056e-20 $X=3.51 $Y=1.03
r127 66 74 4.96191 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=6 $Y=0.95
+ $X2=5.845 $Y2=0.95
r128 65 74 10.404 $w=3.58e-07 $l=3.25e-07 $layer=LI1_cond $X=5.52 $Y=0.95
+ $X2=5.845 $Y2=0.95
r129 65 81 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=5.52 $Y=0.95
+ $X2=5.15 $Y2=0.95
r130 64 81 4.83878 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=0.975
+ $X2=5.15 $Y2=0.975
r131 64 79 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=0.975
+ $X2=4.82 $Y2=0.975
r132 63 66 5.76222 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=6.18 $Y=0.95 $X2=6
+ $Y2=0.95
r133 60 79 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=3.66 $Y=1.095
+ $X2=4.82 $Y2=1.095
r134 54 56 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.565 $Y=0.86
+ $X2=2.565 $Y2=1.03
r135 47 63 8.02311 $w=3.6e-07 $l=2.18403e-07 $layer=LI1_cond $X=6.265 $Y=1.13
+ $X2=6.18 $Y2=0.95
r136 47 48 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.265 $Y=1.13
+ $X2=6.265 $Y2=1.95
r137 46 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.845 $Y=2.035
+ $X2=3.68 $Y2=2.035
r138 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.18 $Y=2.035
+ $X2=6.265 $Y2=1.95
r139 45 46 152.337 $w=1.68e-07 $l=2.335e-06 $layer=LI1_cond $X=6.18 $Y=2.035
+ $X2=3.845 $Y2=2.035
r140 40 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=2.035
+ $X2=2.68 $Y2=2.035
r141 39 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=2.035
+ $X2=3.68 $Y2=2.035
r142 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.515 $Y=2.035
+ $X2=2.845 $Y2=2.035
r143 36 56 1.29116 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=1.03
+ $X2=2.565 $Y2=1.03
r144 36 38 29.3873 $w=2.98e-07 $l=7.65e-07 $layer=LI1_cond $X=2.73 $Y=1.03
+ $X2=3.495 $Y2=1.03
r145 35 60 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.51 $Y=1.03
+ $X2=3.66 $Y2=1.03
r146 35 38 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=3.51 $Y=1.03
+ $X2=3.495 $Y2=1.03
r147 32 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.035
+ $X2=1.68 $Y2=2.035
r148 31 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=2.035
+ $X2=2.68 $Y2=2.035
r149 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.515 $Y=2.035
+ $X2=1.845 $Y2=2.035
r150 28 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r151 27 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=1.68 $Y2=2.035
r152 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=0.945 $Y2=2.035
r153 8 62 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=3.48
+ $Y=1.84 $X2=3.68 $Y2=2.115
r154 7 59 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=1.84 $X2=2.68 $Y2=2.115
r155 6 52 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.115
r156 5 50 300 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.78 $Y2=2.115
r157 4 74 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.37 $X2=5.845 $Y2=0.95
r158 3 64 182 $w=1.7e-07 $l=6.76905e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.37 $X2=4.985 $Y2=0.95
r159 2 38 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.355
+ $Y=0.37 $X2=3.495 $Y2=0.965
r160 1 54 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.37 $X2=2.565 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 50 51 53 54 56 57 58 79 85 86 89
r131 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r132 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r133 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r134 83 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.935 $Y=3.33
+ $X2=9.77 $Y2=3.33
r135 83 85 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.935 $Y=3.33
+ $X2=10.32 $Y2=3.33
r136 82 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r137 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r138 79 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.77 $Y2=3.33
r139 79 81 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.36 $Y2=3.33
r140 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r142 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r143 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r144 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r145 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r146 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r147 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r148 65 66 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r149 62 66 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r150 61 65 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 61 62 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r152 58 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r153 58 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 56 77 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.605 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.605 $Y=3.33
+ $X2=8.77 $Y2=3.33
r156 55 81 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.935 $Y=3.33
+ $X2=9.36 $Y2=3.33
r157 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.935 $Y=3.33
+ $X2=8.77 $Y2=3.33
r158 53 74 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=3.33
+ $X2=7.44 $Y2=3.33
r159 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=3.33
+ $X2=7.77 $Y2=3.33
r160 52 77 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.935 $Y=3.33
+ $X2=8.4 $Y2=3.33
r161 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.935 $Y=3.33
+ $X2=7.77 $Y2=3.33
r162 50 71 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.605 $Y=3.33
+ $X2=6.48 $Y2=3.33
r163 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=3.33
+ $X2=6.77 $Y2=3.33
r164 49 74 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=6.935 $Y=3.33
+ $X2=7.44 $Y2=3.33
r165 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.935 $Y=3.33
+ $X2=6.77 $Y2=3.33
r166 47 68 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.52 $Y2=3.33
r167 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.77 $Y2=3.33
r168 46 71 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.935 $Y=3.33
+ $X2=6.48 $Y2=3.33
r169 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.935 $Y=3.33
+ $X2=5.77 $Y2=3.33
r170 44 65 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.56 $Y2=3.33
r171 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.77 $Y2=3.33
r172 43 68 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=5.52 $Y2=3.33
r173 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=4.77 $Y2=3.33
r174 39 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.77 $Y=3.245
+ $X2=9.77 $Y2=3.33
r175 39 41 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=9.77 $Y=3.245
+ $X2=9.77 $Y2=2.455
r176 35 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.77 $Y=3.245
+ $X2=8.77 $Y2=3.33
r177 35 37 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=8.77 $Y=3.245
+ $X2=8.77 $Y2=2.455
r178 31 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=3.245
+ $X2=7.77 $Y2=3.33
r179 31 33 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=7.77 $Y=3.245
+ $X2=7.77 $Y2=2.455
r180 27 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.77 $Y=3.245
+ $X2=6.77 $Y2=3.33
r181 27 29 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=6.77 $Y=3.245
+ $X2=6.77 $Y2=2.805
r182 23 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.77 $Y=3.245
+ $X2=5.77 $Y2=3.33
r183 23 25 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=5.77 $Y=3.245
+ $X2=5.77 $Y2=2.805
r184 19 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=3.33
r185 19 21 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=2.805
r186 6 41 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=9.57
+ $Y=1.84 $X2=9.77 $Y2=2.455
r187 5 37 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=8.57
+ $Y=1.84 $X2=8.77 $Y2=2.455
r188 4 33 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=7.57
+ $Y=1.84 $X2=7.77 $Y2=2.455
r189 3 29 600 $w=1.7e-07 $l=1.05573e-06 $layer=licon1_PDIFF $count=1 $X=6.58
+ $Y=1.84 $X2=6.77 $Y2=2.805
r190 2 25 600 $w=1.7e-07 $l=1.06029e-06 $layer=licon1_PDIFF $count=1 $X=5.57
+ $Y=1.84 $X2=5.77 $Y2=2.805
r191 1 21 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=4.62
+ $Y=1.84 $X2=4.77 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%A_27_74# 1 2 3 4 5 18 20 21 24 26 32 33 34
+ 36 37 42
c74 32 0 8.60869e-20 $X=2.9 $Y=0.34
r75 42 45 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.925 $Y=0.34
+ $X2=3.925 $Y2=0.53
r76 37 40 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.065 $Y=0.34
+ $X2=3.065 $Y2=0.53
r77 35 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=0.34
+ $X2=3.065 $Y2=0.34
r78 34 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0.34
+ $X2=3.925 $Y2=0.34
r79 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.76 $Y=0.34
+ $X2=3.23 $Y2=0.34
r80 32 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=0.34
+ $X2=3.065 $Y2=0.34
r81 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.9 $Y=0.34 $X2=2.22
+ $Y2=0.34
r82 29 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.135 $Y=1.01
+ $X2=2.135 $Y2=0.515
r83 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=0.425
+ $X2=2.22 $Y2=0.34
r84 28 31 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.135 $Y=0.425
+ $X2=2.135 $Y2=0.515
r85 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=1.095
+ $X2=1.21 $Y2=1.095
r86 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=1.095
+ $X2=2.135 $Y2=1.01
r87 26 27 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.05 $Y=1.095
+ $X2=1.295 $Y2=1.095
r88 22 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=1.01 $X2=1.21
+ $Y2=1.095
r89 22 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.21 $Y=1.01
+ $X2=1.21 $Y2=0.515
r90 20 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=1.21 $Y2=1.095
r91 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=0.445 $Y2=1.095
r92 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r93 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r94 5 45 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.37 $X2=3.925 $Y2=0.53
r95 4 40 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.37 $X2=3.065 $Y2=0.53
r96 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.995
+ $Y=0.37 $X2=2.135 $Y2=0.515
r97 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r98 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 53 58 64 67 70 73 77
r112 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r113 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r114 70 71 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r115 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r116 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r117 62 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r118 62 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r119 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r120 59 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.585 $Y=0 $X2=9.42
+ $Y2=0
r121 59 61 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.585 $Y=0
+ $X2=9.84 $Y2=0
r122 58 76 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.337 $Y2=0
r123 58 61 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.84 $Y2=0
r124 57 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r125 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r126 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r127 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=0 $X2=8.56
+ $Y2=0
r128 54 56 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.725 $Y=0
+ $X2=8.88 $Y2=0
r129 53 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=0 $X2=9.42
+ $Y2=0
r130 53 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.255 $Y=0
+ $X2=8.88 $Y2=0
r131 52 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r132 51 52 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r133 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.64
+ $Y2=0
r134 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=2.16 $Y2=0
r135 48 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.395 $Y=0 $X2=8.56
+ $Y2=0
r136 48 51 406.775 $w=1.68e-07 $l=6.235e-06 $layer=LI1_cond $X=8.395 $Y=0
+ $X2=2.16 $Y2=0
r137 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r138 47 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r139 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r140 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r141 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r142 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.64
+ $Y2=0
r143 43 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r144 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r146 38 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r147 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r148 36 71 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=8.4
+ $Y2=0
r149 36 52 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=2.16 $Y2=0
r150 32 76 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.337 $Y2=0
r151 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0.515
r152 28 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.42 $Y=0.085
+ $X2=9.42 $Y2=0
r153 28 30 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=9.42 $Y=0.085
+ $X2=9.42 $Y2=0.595
r154 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.56 $Y=0.085
+ $X2=8.56 $Y2=0
r155 24 26 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=8.56 $Y=0.085
+ $X2=8.56 $Y2=0.595
r156 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0
r157 20 22 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0.595
r158 16 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r159 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.595
r160 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.14
+ $Y=0.37 $X2=10.28 $Y2=0.515
r161 4 30 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=9.28
+ $Y=0.37 $X2=9.42 $Y2=0.595
r162 3 26 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=8.415
+ $Y=0.37 $X2=8.56 $Y2=0.595
r163 2 22 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.595
r164 1 18 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%A_868_74# 1 2 3 4 5 24 30 31
r40 30 31 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8 $Y=0.515
+ $X2=7.835 $Y2=0.515
r41 24 27 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.485 $Y=0.475
+ $X2=4.485 $Y2=0.595
r42 23 31 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=7.135 $Y=0.475
+ $X2=7.835 $Y2=0.475
r43 21 23 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=6.275 $Y=0.475
+ $X2=7.135 $Y2=0.475
r44 19 21 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=5.415 $Y=0.475
+ $X2=6.275 $Y2=0.475
r45 17 24 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=4.65 $Y=0.475
+ $X2=4.485 $Y2=0.475
r46 17 19 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=4.65 $Y=0.475
+ $X2=5.415 $Y2=0.475
r47 5 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.86
+ $Y=0.37 $X2=8 $Y2=0.515
r48 4 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.995
+ $Y=0.37 $X2=7.135 $Y2=0.515
r49 3 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.135
+ $Y=0.37 $X2=6.275 $Y2=0.515
r50 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.275
+ $Y=0.37 $X2=5.415 $Y2=0.515
r51 1 27 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.37 $X2=4.485 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_4%A_1313_74# 1 2 3 4 15 19 21 25 30 32 33 34
r57 32 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.57 $Y=1.015
+ $X2=7.735 $Y2=1.015
r58 30 32 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=6.87 $Y=1.015 $X2=7.57
+ $Y2=1.015
r59 28 30 5.11015 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.705 $Y=0.975
+ $X2=6.87 $Y2=0.975
r60 23 25 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.85 $Y=1.01
+ $X2=9.85 $Y2=0.515
r61 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.075 $Y=1.095
+ $X2=8.99 $Y2=1.095
r62 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.765 $Y=1.095
+ $X2=9.85 $Y2=1.01
r63 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.765 $Y=1.095
+ $X2=9.075 $Y2=1.095
r64 17 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=1.01 $X2=8.99
+ $Y2=1.095
r65 17 19 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.99 $Y=1.01
+ $X2=8.99 $Y2=0.515
r66 15 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=1.095
+ $X2=8.99 $Y2=1.095
r67 15 33 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=8.905 $Y=1.095
+ $X2=7.735 $Y2=1.095
r68 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.71
+ $Y=0.37 $X2=9.85 $Y2=0.515
r69 3 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.85
+ $Y=0.37 $X2=8.99 $Y2=0.515
r70 2 32 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=7.43
+ $Y=0.37 $X2=7.57 $Y2=0.95
r71 1 28 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.37 $X2=6.705 $Y2=0.95
.ends

