* File: sky130_fd_sc_hs__o21ai_1.spice
* Created: Tue Sep  1 20:14:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o21ai_1.pex.spice"
.subckt sky130_fd_sc_hs__o21ai_1  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_27_74#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3361 AS=0.2109 PD=1.68 PS=2.05 NRD=64.728 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1001 N_A_27_74#_M1001_d N_A2_M1001_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3361 PD=1.02 PS=1.68 NRD=0 NRS=64.728 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_27_74#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1005 A_162_368# N_A1_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.4648 PD=1.39 PS=3.07 NRD=14.0658 NRS=8.7862 M=1 R=7.46667 SA=75000.3
+ SB=75001.3 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_A2_M1000_g A_162_368# VPB PSHORT L=0.15 W=1.12 AD=0.2828
+ AS=0.1512 PD=1.625 PS=1.39 NRD=1.7533 NRS=14.0658 M=1 R=7.46667 SA=75000.8
+ SB=75000.9 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_Y_M1000_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2828 PD=2.83 PS=1.625 NRD=1.7533 NRS=37.8043 M=1 R=7.46667
+ SA=75001.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_hs__o21ai_1.pxi.spice"
*
.ends
*
*
