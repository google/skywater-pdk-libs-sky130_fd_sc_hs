* File: sky130_fd_sc_hs__and4b_1.pxi.spice
* Created: Thu Aug 27 20:33:24 2020
* 
x_PM_SKY130_FD_SC_HS__AND4B_1%A_N N_A_N_M1010_g N_A_N_c_85_n N_A_N_M1009_g
+ N_A_N_c_82_n A_N N_A_N_c_83_n N_A_N_c_84_n PM_SKY130_FD_SC_HS__AND4B_1%A_N
x_PM_SKY130_FD_SC_HS__AND4B_1%A_27_74# N_A_27_74#_M1010_s N_A_27_74#_M1009_s
+ N_A_27_74#_c_119_n N_A_27_74#_M1008_g N_A_27_74#_c_120_n N_A_27_74#_c_121_n
+ N_A_27_74#_c_122_n N_A_27_74#_c_123_n N_A_27_74#_M1006_g N_A_27_74#_c_124_n
+ N_A_27_74#_c_130_n N_A_27_74#_c_125_n N_A_27_74#_c_126_n N_A_27_74#_c_131_n
+ N_A_27_74#_c_132_n N_A_27_74#_c_127_n N_A_27_74#_c_133_n N_A_27_74#_c_128_n
+ PM_SKY130_FD_SC_HS__AND4B_1%A_27_74#
x_PM_SKY130_FD_SC_HS__AND4B_1%B N_B_c_204_n N_B_M1005_g N_B_M1003_g N_B_c_201_n
+ N_B_c_202_n B B PM_SKY130_FD_SC_HS__AND4B_1%B
x_PM_SKY130_FD_SC_HS__AND4B_1%C N_C_M1011_g N_C_c_238_n N_C_c_243_n N_C_M1001_g
+ N_C_c_239_n C C N_C_c_240_n N_C_c_241_n PM_SKY130_FD_SC_HS__AND4B_1%C
x_PM_SKY130_FD_SC_HS__AND4B_1%D N_D_c_284_n N_D_M1002_g N_D_M1000_g D
+ PM_SKY130_FD_SC_HS__AND4B_1%D
x_PM_SKY130_FD_SC_HS__AND4B_1%A_226_424# N_A_226_424#_M1006_s
+ N_A_226_424#_M1008_d N_A_226_424#_M1001_d N_A_226_424#_c_321_n
+ N_A_226_424#_M1004_g N_A_226_424#_c_322_n N_A_226_424#_M1007_g
+ N_A_226_424#_c_323_n N_A_226_424#_c_324_n N_A_226_424#_c_325_n
+ N_A_226_424#_c_326_n N_A_226_424#_c_327_n N_A_226_424#_c_331_n
+ N_A_226_424#_c_333_n N_A_226_424#_c_367_n N_A_226_424#_c_354_n
+ N_A_226_424#_c_332_n PM_SKY130_FD_SC_HS__AND4B_1%A_226_424#
x_PM_SKY130_FD_SC_HS__AND4B_1%VPWR N_VPWR_M1009_d N_VPWR_M1005_d N_VPWR_M1002_d
+ N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n VPWR
+ N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_419_n N_VPWR_c_427_n N_VPWR_c_428_n
+ N_VPWR_c_429_n PM_SKY130_FD_SC_HS__AND4B_1%VPWR
x_PM_SKY130_FD_SC_HS__AND4B_1%X N_X_M1007_d N_X_M1004_d N_X_c_466_n N_X_c_467_n
+ X X X X N_X_c_468_n PM_SKY130_FD_SC_HS__AND4B_1%X
x_PM_SKY130_FD_SC_HS__AND4B_1%VGND N_VGND_M1010_d N_VGND_M1000_d N_VGND_c_491_n
+ N_VGND_c_492_n VGND N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n
+ N_VGND_c_496_n N_VGND_c_497_n N_VGND_c_498_n PM_SKY130_FD_SC_HS__AND4B_1%VGND
cc_1 VNB N_A_N_M1010_g 0.0371391f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_A_N_c_82_n 0.0249613f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.695
cc_3 VNB N_A_N_c_83_n 0.0184956f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_4 VNB N_A_N_c_84_n 0.0229758f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_5 VNB N_A_27_74#_c_119_n 0.0174436f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_6 VNB N_A_27_74#_c_120_n 0.0668854f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_27_74#_c_121_n 0.0305639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_122_n 0.0108824f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_9 VNB N_A_27_74#_c_123_n 0.0132493f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_10 VNB N_A_27_74#_c_124_n 0.0214334f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.525
cc_11 VNB N_A_27_74#_c_125_n 0.0105312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_126_n 0.00992961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_127_n 0.0108784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_128_n 0.00226763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_M1003_g 0.0301282f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_16 VNB N_B_c_201_n 0.0158533f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_17 VNB N_B_c_202_n 0.0334807f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.19
cc_18 VNB B 0.00854044f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_C_M1011_g 0.00933542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_c_238_n 0.0196984f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_21 VNB N_C_c_239_n 0.0158129f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_C_c_240_n 0.0412509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_241_n 0.025844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_D_c_284_n 0.0269821f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.19
cc_25 VNB N_D_M1000_g 0.0298855f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_26 VNB D 0.00251027f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_27 VNB N_A_226_424#_c_321_n 0.0279356f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.695
cc_28 VNB N_A_226_424#_c_322_n 0.0215792f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_29 VNB N_A_226_424#_c_323_n 0.00846748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_226_424#_c_324_n 0.00939658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_226_424#_c_325_n 0.0105635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_226_424#_c_326_n 0.00482938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_226_424#_c_327_n 0.0214217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_419_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_466_n 0.0240518f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.19
cc_36 VNB N_X_c_467_n 0.00694384f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_37 VNB N_X_c_468_n 0.0219872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_491_n 0.0175884f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.19
cc_39 VNB N_VGND_c_492_n 0.0190854f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_40 VNB N_VGND_c_493_n 0.0181399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_494_n 0.0705391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_495_n 0.019578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_496_n 0.293095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_497_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_498_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_A_N_c_85_n 0.0202931f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_47 VPB N_A_N_c_82_n 0.0364599f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.695
cc_48 VPB N_A_N_c_84_n 0.0103985f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.355
cc_49 VPB N_A_27_74#_c_119_n 0.0473337f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_50 VPB N_A_27_74#_c_130_n 0.0323583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_27_74#_c_131_n 0.0074636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_27_74#_c_132_n 0.00998527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_74#_c_133_n 0.0032226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_74#_c_128_n 0.00358177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_B_c_204_n 0.0200481f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.19
cc_56 VPB N_B_c_201_n 0.00910323f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.355
cc_57 VPB N_B_c_202_n 0.0153875f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.19
cc_58 VPB B 4.81172e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_59 VPB N_C_c_238_n 7.66471e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_60 VPB N_C_c_243_n 0.0273103f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_61 VPB N_D_c_284_n 0.0374717f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.19
cc_62 VPB D 0.00257344f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.355
cc_63 VPB N_A_226_424#_c_321_n 0.034579f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.695
cc_64 VPB N_A_226_424#_c_326_n 0.00181129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_226_424#_c_327_n 0.00422694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_226_424#_c_331_n 0.00289255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_226_424#_c_332_n 0.00870398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_420_n 0.009836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_421_n 0.0157802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_422_n 0.0207378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_423_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_424_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_425_n 0.0202291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_419_n 0.0789208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_427_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_428_n 0.0220529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_429_n 0.0277939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB X 0.00694384f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.355
cc_79 VPB X 0.0403408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_X_c_468_n 0.00914129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 N_A_N_c_85_n N_A_27_74#_c_119_n 0.0230192f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_82 N_A_N_c_82_n N_A_27_74#_c_119_n 0.0160755f $X=0.43 $Y=1.695 $X2=0 $Y2=0
cc_83 N_A_N_c_84_n N_A_27_74#_c_119_n 3.08399e-19 $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_84 N_A_N_c_83_n N_A_27_74#_c_120_n 0.00596009f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_85 N_A_N_M1010_g N_A_27_74#_c_122_n 0.0114901f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_86 N_A_N_M1010_g N_A_27_74#_c_124_n 0.00226722f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_87 N_A_N_c_85_n N_A_27_74#_c_130_n 0.0129585f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_88 N_A_N_M1010_g N_A_27_74#_c_125_n 0.0140234f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_89 N_A_N_c_83_n N_A_27_74#_c_125_n 0.00104829f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_90 N_A_N_c_84_n N_A_27_74#_c_125_n 0.0144955f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_91 N_A_N_c_83_n N_A_27_74#_c_126_n 0.00375152f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_92 N_A_N_c_84_n N_A_27_74#_c_126_n 0.0254263f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_93 N_A_N_c_85_n N_A_27_74#_c_131_n 0.00997674f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_94 N_A_N_c_82_n N_A_27_74#_c_131_n 0.00268084f $X=0.43 $Y=1.695 $X2=0 $Y2=0
cc_95 N_A_N_c_84_n N_A_27_74#_c_131_n 0.0113214f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_96 N_A_N_c_85_n N_A_27_74#_c_132_n 0.00169587f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_97 N_A_N_c_82_n N_A_27_74#_c_132_n 0.0051831f $X=0.43 $Y=1.695 $X2=0 $Y2=0
cc_98 N_A_N_c_84_n N_A_27_74#_c_132_n 0.0288658f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_99 N_A_N_M1010_g N_A_27_74#_c_127_n 0.00374114f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_100 N_A_N_c_83_n N_A_27_74#_c_127_n 0.0013621f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_101 N_A_N_c_84_n N_A_27_74#_c_127_n 0.0266416f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_102 N_A_N_c_82_n N_A_27_74#_c_133_n 0.00321029f $X=0.43 $Y=1.695 $X2=0 $Y2=0
cc_103 N_A_N_c_82_n N_A_27_74#_c_128_n 0.00172483f $X=0.43 $Y=1.695 $X2=0 $Y2=0
cc_104 N_A_N_c_84_n N_A_27_74#_c_128_n 0.0248669f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_105 N_A_N_c_85_n N_A_226_424#_c_333_n 5.87414e-19 $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_106 N_A_N_c_85_n N_VPWR_c_420_n 0.00689824f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_107 N_A_N_c_85_n N_VPWR_c_424_n 0.00445602f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_108 N_A_N_c_85_n N_VPWR_c_419_n 0.00861319f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_109 N_A_N_M1010_g N_VGND_c_491_n 0.00527104f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_110 N_A_N_M1010_g N_VGND_c_493_n 0.00461464f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_111 N_A_N_M1010_g N_VGND_c_496_n 0.00473629f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_112 N_A_27_74#_c_119_n N_B_c_204_n 0.0250912f $X=1.055 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_27_74#_c_123_n N_B_M1003_g 0.0314813f $X=1.69 $Y=0.545 $X2=0 $Y2=0
cc_114 N_A_27_74#_c_119_n N_B_c_201_n 0.0202716f $X=1.055 $Y=2.045 $X2=0 $Y2=0
cc_115 N_A_27_74#_c_123_n N_B_c_201_n 0.00834499f $X=1.69 $Y=0.545 $X2=0 $Y2=0
cc_116 N_A_27_74#_c_128_n N_B_c_201_n 0.00110467f $X=1.09 $Y=1.715 $X2=0 $Y2=0
cc_117 N_A_27_74#_c_119_n B 0.00114193f $X=1.055 $Y=2.045 $X2=0 $Y2=0
cc_118 N_A_27_74#_c_123_n B 0.00104663f $X=1.69 $Y=0.545 $X2=0 $Y2=0
cc_119 N_A_27_74#_c_133_n B 0.00232826f $X=0.86 $Y=2.03 $X2=0 $Y2=0
cc_120 N_A_27_74#_c_128_n B 0.0170835f $X=1.09 $Y=1.715 $X2=0 $Y2=0
cc_121 N_A_27_74#_c_121_n N_C_c_240_n 0.00170036f $X=1.615 $Y=0.47 $X2=0 $Y2=0
cc_122 N_A_27_74#_c_121_n N_C_c_241_n 0.00647686f $X=1.615 $Y=0.47 $X2=0 $Y2=0
cc_123 N_A_27_74#_c_120_n N_A_226_424#_c_323_n 0.0099514f $X=1.18 $Y=1.55 $X2=0
+ $Y2=0
cc_124 N_A_27_74#_c_121_n N_A_226_424#_c_323_n 0.0052648f $X=1.615 $Y=0.47 $X2=0
+ $Y2=0
cc_125 N_A_27_74#_c_123_n N_A_226_424#_c_323_n 0.0119422f $X=1.69 $Y=0.545 $X2=0
+ $Y2=0
cc_126 N_A_27_74#_c_125_n N_A_226_424#_c_323_n 0.0088137f $X=0.775 $Y=0.935
+ $X2=0 $Y2=0
cc_127 N_A_27_74#_c_127_n N_A_226_424#_c_323_n 0.00880168f $X=0.86 $Y=1.55 $X2=0
+ $Y2=0
cc_128 N_A_27_74#_c_123_n N_A_226_424#_c_324_n 0.0102279f $X=1.69 $Y=0.545 $X2=0
+ $Y2=0
cc_129 N_A_27_74#_c_120_n N_A_226_424#_c_325_n 0.00218369f $X=1.18 $Y=1.55 $X2=0
+ $Y2=0
cc_130 N_A_27_74#_c_123_n N_A_226_424#_c_325_n 0.00196337f $X=1.69 $Y=0.545
+ $X2=0 $Y2=0
cc_131 N_A_27_74#_c_127_n N_A_226_424#_c_325_n 0.00841426f $X=0.86 $Y=1.55 $X2=0
+ $Y2=0
cc_132 N_A_27_74#_c_119_n N_A_226_424#_c_333_n 0.00838744f $X=1.055 $Y=2.045
+ $X2=0 $Y2=0
cc_133 N_A_27_74#_c_130_n N_A_226_424#_c_333_n 0.00425759f $X=0.28 $Y=2.265
+ $X2=0 $Y2=0
cc_134 N_A_27_74#_c_128_n N_A_226_424#_c_333_n 0.00629839f $X=1.09 $Y=1.715
+ $X2=0 $Y2=0
cc_135 N_A_27_74#_c_131_n N_VPWR_M1009_d 0.00370145f $X=0.775 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_27_74#_c_119_n N_VPWR_c_420_n 0.00727882f $X=1.055 $Y=2.045 $X2=0
+ $Y2=0
cc_137 N_A_27_74#_c_130_n N_VPWR_c_420_n 0.0236791f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_138 N_A_27_74#_c_131_n N_VPWR_c_420_n 0.023834f $X=0.775 $Y=2.115 $X2=0 $Y2=0
cc_139 N_A_27_74#_c_130_n N_VPWR_c_424_n 0.0145938f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_140 N_A_27_74#_c_119_n N_VPWR_c_419_n 0.00909941f $X=1.055 $Y=2.045 $X2=0
+ $Y2=0
cc_141 N_A_27_74#_c_130_n N_VPWR_c_419_n 0.0120466f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_142 N_A_27_74#_c_119_n N_VPWR_c_428_n 0.00461464f $X=1.055 $Y=2.045 $X2=0
+ $Y2=0
cc_143 N_A_27_74#_c_119_n N_VPWR_c_429_n 0.00252936f $X=1.055 $Y=2.045 $X2=0
+ $Y2=0
cc_144 N_A_27_74#_c_125_n N_VGND_M1010_d 0.0025118f $X=0.775 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_27_74#_c_122_n N_VGND_c_491_n 0.0059979f $X=1.255 $Y=0.47 $X2=0 $Y2=0
cc_146 N_A_27_74#_c_124_n N_VGND_c_491_n 0.00155433f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_147 N_A_27_74#_c_125_n N_VGND_c_491_n 0.0206247f $X=0.775 $Y=0.935 $X2=0
+ $Y2=0
cc_148 N_A_27_74#_c_124_n N_VGND_c_493_n 0.0128369f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_149 N_A_27_74#_c_122_n N_VGND_c_494_n 0.017157f $X=1.255 $Y=0.47 $X2=0 $Y2=0
cc_150 N_A_27_74#_c_122_n N_VGND_c_496_n 0.0206598f $X=1.255 $Y=0.47 $X2=0 $Y2=0
cc_151 N_A_27_74#_c_124_n N_VGND_c_496_n 0.0106314f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_152 N_A_27_74#_c_125_n N_VGND_c_496_n 0.00853677f $X=0.775 $Y=0.935 $X2=0
+ $Y2=0
cc_153 N_B_M1003_g N_C_c_238_n 0.00693254f $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_154 B N_C_c_238_n 0.00297314f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_155 N_B_c_202_n N_C_c_243_n 0.00693254f $X=2.09 $Y=1.795 $X2=0 $Y2=0
cc_156 N_B_M1003_g N_C_c_240_n 0.0564627f $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_157 N_B_M1003_g N_C_c_241_n 0.0101643f $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_158 N_B_M1003_g N_A_226_424#_c_323_n 0.00265403f $X=2.165 $Y=1.015 $X2=0
+ $Y2=0
cc_159 N_B_M1003_g N_A_226_424#_c_324_n 0.0122201f $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_160 N_B_c_202_n N_A_226_424#_c_324_n 0.00185324f $X=2.09 $Y=1.795 $X2=0 $Y2=0
cc_161 B N_A_226_424#_c_324_n 0.0495197f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_162 N_B_c_201_n N_A_226_424#_c_325_n 0.00341415f $X=1.675 $Y=1.795 $X2=0
+ $Y2=0
cc_163 B N_A_226_424#_c_325_n 0.00662497f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_164 N_B_M1003_g N_A_226_424#_c_326_n 0.00133983f $X=2.165 $Y=1.015 $X2=0
+ $Y2=0
cc_165 B N_A_226_424#_c_326_n 0.0206392f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_166 N_B_c_204_n N_A_226_424#_c_354_n 0.0215994f $X=1.585 $Y=2.045 $X2=0 $Y2=0
cc_167 N_B_c_202_n N_A_226_424#_c_354_n 0.0131963f $X=2.09 $Y=1.795 $X2=0 $Y2=0
cc_168 B N_A_226_424#_c_354_n 0.0520232f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_169 N_B_c_204_n N_VPWR_c_419_n 0.00813866f $X=1.585 $Y=2.045 $X2=0 $Y2=0
cc_170 N_B_c_204_n N_VPWR_c_428_n 0.00413917f $X=1.585 $Y=2.045 $X2=0 $Y2=0
cc_171 N_B_c_204_n N_VPWR_c_429_n 0.0170483f $X=1.585 $Y=2.045 $X2=0 $Y2=0
cc_172 N_B_M1003_g N_VGND_c_494_n 4.64175e-19 $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_173 N_C_c_238_n N_D_c_284_n 0.00581811f $X=2.655 $Y=1.955 $X2=-0.19
+ $Y2=-0.245
cc_174 N_C_c_243_n N_D_c_284_n 0.0207021f $X=2.655 $Y=2.045 $X2=-0.19 $Y2=-0.245
cc_175 N_C_c_239_n N_D_c_284_n 0.017484f $X=2.612 $Y=1.56 $X2=-0.19 $Y2=-0.245
cc_176 N_C_M1011_g N_D_M1000_g 0.0197345f $X=2.555 $Y=1.015 $X2=0 $Y2=0
cc_177 N_C_c_239_n N_D_M1000_g 0.00334362f $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_178 N_C_c_240_n N_D_M1000_g 0.0034753f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_179 N_C_c_241_n N_D_M1000_g 0.00131309f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_180 N_C_c_239_n D 4.09211e-19 $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_181 N_C_c_241_n N_A_226_424#_c_323_n 0.0030474f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_182 N_C_M1011_g N_A_226_424#_c_324_n 0.0110133f $X=2.555 $Y=1.015 $X2=0 $Y2=0
cc_183 N_C_c_241_n N_A_226_424#_c_324_n 0.0149142f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_184 N_C_M1011_g N_A_226_424#_c_326_n 8.15891e-19 $X=2.555 $Y=1.015 $X2=0
+ $Y2=0
cc_185 N_C_c_238_n N_A_226_424#_c_326_n 0.0100704f $X=2.655 $Y=1.955 $X2=0 $Y2=0
cc_186 N_C_c_243_n N_A_226_424#_c_326_n 0.00843863f $X=2.655 $Y=2.045 $X2=0
+ $Y2=0
cc_187 N_C_c_239_n N_A_226_424#_c_326_n 0.00724776f $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_188 N_C_c_240_n N_A_226_424#_c_327_n 2.05086e-19 $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_189 N_C_c_241_n N_A_226_424#_c_327_n 0.00154757f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_190 N_C_c_243_n N_A_226_424#_c_331_n 0.00341623f $X=2.655 $Y=2.045 $X2=0
+ $Y2=0
cc_191 N_C_M1011_g N_A_226_424#_c_367_n 0.00463728f $X=2.555 $Y=1.015 $X2=0
+ $Y2=0
cc_192 N_C_c_240_n N_A_226_424#_c_367_n 5.51222e-19 $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_193 N_C_c_241_n N_A_226_424#_c_367_n 0.00519212f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_194 N_C_c_243_n N_A_226_424#_c_354_n 0.00637947f $X=2.655 $Y=2.045 $X2=0
+ $Y2=0
cc_195 N_C_c_239_n N_A_226_424#_c_354_n 0.00187615f $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_196 N_C_c_243_n N_A_226_424#_c_332_n 0.0145626f $X=2.655 $Y=2.045 $X2=0 $Y2=0
cc_197 N_C_c_243_n N_VPWR_c_422_n 0.00413917f $X=2.655 $Y=2.045 $X2=0 $Y2=0
cc_198 N_C_c_243_n N_VPWR_c_419_n 0.00813626f $X=2.655 $Y=2.045 $X2=0 $Y2=0
cc_199 N_C_c_243_n N_VPWR_c_429_n 0.0120728f $X=2.655 $Y=2.045 $X2=0 $Y2=0
cc_200 N_C_c_240_n N_VGND_c_492_n 0.00126694f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_201 N_C_c_241_n N_VGND_c_492_n 0.0130106f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_202 N_C_c_240_n N_VGND_c_494_n 0.00783549f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_203 N_C_c_241_n N_VGND_c_494_n 0.0514254f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_204 N_C_c_240_n N_VGND_c_496_n 0.011167f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_205 N_C_c_241_n N_VGND_c_496_n 0.0291589f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_206 N_D_c_284_n N_A_226_424#_c_321_n 0.0257962f $X=3.155 $Y=2.045 $X2=0 $Y2=0
cc_207 N_D_M1000_g N_A_226_424#_c_321_n 0.0170787f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_208 D N_A_226_424#_c_321_n 0.00123715f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_209 N_D_M1000_g N_A_226_424#_c_322_n 0.0185769f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_210 N_D_c_284_n N_A_226_424#_c_326_n 0.00585751f $X=3.155 $Y=2.045 $X2=0
+ $Y2=0
cc_211 N_D_M1000_g N_A_226_424#_c_326_n 0.00283662f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_212 D N_A_226_424#_c_326_n 0.0204438f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_213 N_D_c_284_n N_A_226_424#_c_327_n 0.00128789f $X=3.155 $Y=2.045 $X2=0
+ $Y2=0
cc_214 N_D_M1000_g N_A_226_424#_c_327_n 0.021225f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_215 D N_A_226_424#_c_327_n 0.032803f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_216 N_D_c_284_n N_A_226_424#_c_331_n 0.00957895f $X=3.155 $Y=2.045 $X2=0
+ $Y2=0
cc_217 N_D_c_284_n N_A_226_424#_c_332_n 0.0043602f $X=3.155 $Y=2.045 $X2=0 $Y2=0
cc_218 D N_A_226_424#_c_332_n 0.00692482f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_219 N_D_c_284_n N_VPWR_c_421_n 0.012148f $X=3.155 $Y=2.045 $X2=0 $Y2=0
cc_220 N_D_c_284_n N_VPWR_c_422_n 0.00445602f $X=3.155 $Y=2.045 $X2=0 $Y2=0
cc_221 N_D_c_284_n N_VPWR_c_419_n 0.00860522f $X=3.155 $Y=2.045 $X2=0 $Y2=0
cc_222 N_D_c_284_n N_VPWR_c_429_n 6.6728e-19 $X=3.155 $Y=2.045 $X2=0 $Y2=0
cc_223 N_D_M1000_g N_X_c_466_n 7.43364e-19 $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_224 N_D_c_284_n X 8.30284e-19 $X=3.155 $Y=2.045 $X2=0 $Y2=0
cc_225 D X 8.49296e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_226 N_D_c_284_n X 4.02232e-19 $X=3.155 $Y=2.045 $X2=0 $Y2=0
cc_227 N_D_M1000_g N_VGND_c_492_n 0.00462414f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_228 N_D_M1000_g N_VGND_c_494_n 0.00428744f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_229 N_D_M1000_g N_VGND_c_496_n 0.00476395f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_230 N_A_226_424#_c_354_n N_VPWR_M1005_d 0.0290639f $X=2.595 $Y=2.225 $X2=0
+ $Y2=0
cc_231 N_A_226_424#_c_321_n N_VPWR_c_421_n 0.0130989f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_226_424#_c_327_n N_VPWR_c_421_n 0.00555466f $X=3.535 $Y=1.295 $X2=0
+ $Y2=0
cc_233 N_A_226_424#_c_331_n N_VPWR_c_421_n 0.0375649f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_234 N_A_226_424#_c_332_n N_VPWR_c_421_n 0.0156418f $X=2.93 $Y=2.265 $X2=0
+ $Y2=0
cc_235 N_A_226_424#_c_331_n N_VPWR_c_422_n 0.014513f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_236 N_A_226_424#_c_321_n N_VPWR_c_425_n 0.00445602f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A_226_424#_c_321_n N_VPWR_c_419_n 0.00862964f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_226_424#_c_331_n N_VPWR_c_419_n 0.0120152f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_239 N_A_226_424#_c_331_n N_VPWR_c_429_n 0.0194969f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_240 N_A_226_424#_c_354_n N_VPWR_c_429_n 0.0644485f $X=2.595 $Y=2.225 $X2=0
+ $Y2=0
cc_241 N_A_226_424#_c_322_n N_X_c_466_n 0.00609418f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_242 N_A_226_424#_c_322_n N_X_c_467_n 0.00371672f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_243 N_A_226_424#_c_327_n N_X_c_467_n 0.001126f $X=3.535 $Y=1.295 $X2=0 $Y2=0
cc_244 N_A_226_424#_c_321_n X 0.00380226f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_226_424#_c_327_n X 0.00108105f $X=3.535 $Y=1.295 $X2=0 $Y2=0
cc_246 N_A_226_424#_c_321_n X 0.0118888f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_247 N_A_226_424#_c_321_n N_X_c_468_n 0.0117962f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A_226_424#_c_322_n N_X_c_468_n 0.00255066f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_249 N_A_226_424#_c_327_n N_X_c_468_n 0.0309163f $X=3.535 $Y=1.295 $X2=0 $Y2=0
cc_250 N_A_226_424#_c_327_n N_VGND_M1000_d 0.00339782f $X=3.535 $Y=1.295 $X2=0
+ $Y2=0
cc_251 N_A_226_424#_c_323_n N_VGND_c_491_n 0.00343679f $X=1.475 $Y=0.765 $X2=0
+ $Y2=0
cc_252 N_A_226_424#_c_321_n N_VGND_c_492_n 7.86248e-19 $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_253 N_A_226_424#_c_322_n N_VGND_c_492_n 0.00807563f $X=3.825 $Y=1.35 $X2=0
+ $Y2=0
cc_254 N_A_226_424#_c_327_n N_VGND_c_492_n 0.026684f $X=3.535 $Y=1.295 $X2=0
+ $Y2=0
cc_255 N_A_226_424#_c_323_n N_VGND_c_494_n 0.00707634f $X=1.475 $Y=0.765 $X2=0
+ $Y2=0
cc_256 N_A_226_424#_c_322_n N_VGND_c_495_n 0.00467453f $X=3.825 $Y=1.35 $X2=0
+ $Y2=0
cc_257 N_A_226_424#_c_322_n N_VGND_c_496_n 0.00505379f $X=3.825 $Y=1.35 $X2=0
+ $Y2=0
cc_258 N_A_226_424#_c_323_n N_VGND_c_496_n 0.0101843f $X=1.475 $Y=0.765 $X2=0
+ $Y2=0
cc_259 N_A_226_424#_c_324_n A_353_124# 0.00805082f $X=2.595 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_226_424#_c_324_n A_448_139# 0.00237138f $X=2.595 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_261 N_A_226_424#_c_327_n A_526_139# 0.0125125f $X=3.535 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_262 N_A_226_424#_c_367_n A_526_139# 0.00134898f $X=2.68 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_263 N_VPWR_c_421_n X 0.0584082f $X=3.5 $Y=2.265 $X2=0 $Y2=0
cc_264 N_VPWR_c_425_n X 0.0157093f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_265 N_VPWR_c_419_n X 0.0129699f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_266 N_X_c_466_n N_VGND_c_492_n 0.0220013f $X=4.04 $Y=0.645 $X2=0 $Y2=0
cc_267 N_X_c_466_n N_VGND_c_495_n 0.0102463f $X=4.04 $Y=0.645 $X2=0 $Y2=0
cc_268 N_X_c_466_n N_VGND_c_496_n 0.0119585f $X=4.04 $Y=0.645 $X2=0 $Y2=0
