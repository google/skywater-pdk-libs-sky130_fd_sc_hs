* NGSPICE file created from sky130_fd_sc_hs__xnor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xnor3_1 A B C VGND VNB VPB VPWR X
M1000 a_786_100# B VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.0267e+12p ps=7.95e+06u
M1001 VPWR a_81_268# X VPB pshort w=1.12e+06u l=150000u
+  ad=1.2852e+12p pd=9.15e+06u as=3.192e+11p ps=2.81e+06u
M1002 VGND a_81_268# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1003 a_1113_383# B a_371_74# VNB nlowvt w=640000u l=150000u
+  ad=4.096e+11p pd=3.95e+06u as=4.48e+11p ps=3.96e+06u
M1004 a_897_54# B a_371_74# VPB pshort w=840000u l=150000u
+  ad=7.3745e+11p pd=5.65e+06u as=6.14e+11p ps=4.91e+06u
M1005 a_371_74# a_232_162# a_81_268# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=4.1795e+11p ps=2.85e+06u
M1006 VPWR A a_897_54# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_1113_383# a_897_54# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_363_394# a_232_162# a_81_268# VNB nlowvt w=640000u l=150000u
+  ad=4.271e+11p pd=3.96e+06u as=2.24e+11p ps=1.98e+06u
M1009 a_786_100# B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1010 a_371_74# a_786_100# a_897_54# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.95425e+11p ps=4.74e+06u
M1011 a_81_268# C a_371_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_232_162# C VPWR VPB pshort w=640000u l=150000u
+  ad=1.888e+11p pd=1.87e+06u as=0p ps=0u
M1013 a_232_162# C VGND VNB nlowvt w=420000u l=150000u
+  ad=1.575e+11p pd=1.59e+06u as=0p ps=0u
M1014 a_81_268# C a_363_394# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=5.532e+11p ps=4.72e+06u
M1015 a_897_54# B a_363_394# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_363_394# a_786_100# a_897_54# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1113_383# B a_363_394# VPB pshort w=640000u l=150000u
+  ad=4.92e+11p pd=4.48e+06u as=0p ps=0u
M1018 a_1113_383# a_897_54# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_371_74# a_786_100# a_1113_383# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A a_897_54# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_363_394# a_786_100# a_1113_383# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

