* File: sky130_fd_sc_hs__dlclkp_2.spice
* Created: Tue Sep  1 20:01:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlclkp_2.pex.spice"
.subckt sky130_fd_sc_hs__dlclkp_2  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_A_83_244#_M1020_g N_A_27_74#_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.224467 AS=0.2109 PD=1.45319 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1014 A_267_74# N_GATE_M1014_g N_VGND_M1020_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.194133 PD=0.88 PS=1.25681 NRD=12.18 NRS=62.808 M=1 R=4.26667
+ SA=75001 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_83_244#_M1013_d N_A_315_48#_M1013_g A_267_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.184091 AS=0.0768 PD=1.49132 PS=0.88 NRD=22.488 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1006 A_494_118# N_A_315_338#_M1006_g N_A_83_244#_M1013_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0774375 AS=0.120809 PD=0.85 PS=0.978679 NRD=36.96 NRS=55.704 M=1
+ R=2.8 SA=75002.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_27_74#_M1010_g A_494_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.125529 AS=0.0774375 PD=0.99569 PS=0.85 NRD=0 NRS=36.96 M=1 R=2.8 SA=75002
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1011 N_A_315_338#_M1011_d N_A_315_48#_M1011_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.221171 PD=2.05 PS=1.75431 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_CLK_M1015_g N_A_315_48#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1019 A_1044_119# N_CLK_M1019_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0777 AS=0.1295 PD=0.95 PS=1.09 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_1041_387#_M1018_d N_A_27_74#_M1018_g A_1044_119# VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.0777 PD=2.05 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_GCLK_M1001_d N_A_1041_387#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.21835 PD=1.02 PS=2.21 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_GCLK_M1001_d N_A_1041_387#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VPWR_M1012_d N_A_83_244#_M1012_g N_A_27_74#_M1012_s VPB PSHORT L=0.15
+ W=1.12 AD=0.328498 AS=0.3304 PD=1.80679 PS=2.83 NRD=28.1316 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75002 A=0.168 P=2.54 MULT=1
MM1000 A_264_392# N_GATE_M1000_g N_VPWR_M1012_d VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.293302 PD=1.27 PS=1.61321 NRD=15.7403 NRS=29.55 M=1 R=6.66667 SA=75001
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1004 N_A_83_244#_M1004_d N_A_315_338#_M1004_g A_264_392# VPB PSHORT L=0.15 W=1
+ AD=0.300493 AS=0.135 PD=2.32394 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.4 SB=75001 A=0.15 P=2.3 MULT=1
MM1007 A_508_508# N_A_315_48#_M1007_g N_A_83_244#_M1004_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.126207 PD=0.69 PS=0.976056 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75002.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_27_74#_M1021_g A_508_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0567 PD=0.933333 PS=0.69 NRD=53.9386 NRS=37.5088 M=1 R=2.8
+ SA=75002.6 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1016 N_A_315_338#_M1016_d N_A_315_48#_M1016_g N_VPWR_M1021_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.231 PD=2.27 PS=1.86667 NRD=2.3443 NRS=38.6908 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_CLK_M1002_g N_A_315_48#_M1002_s VPB PSHORT L=0.15 W=0.84
+ AD=0.155491 AS=0.2646 PD=1.23717 PS=2.31 NRD=9.3772 NRS=7.0329 M=1 R=5.6
+ SA=75000.2 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1017 N_A_1041_387#_M1017_d N_CLK_M1017_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1
+ AD=0.1625 AS=0.185109 PD=1.325 PS=1.47283 NRD=6.8753 NRS=6.8753 M=1 R=6.66667
+ SA=75000.7 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_27_74#_M1009_g N_A_1041_387#_M1017_d VPB PSHORT L=0.15
+ W=1 AD=0.473255 AS=0.1625 PD=1.9717 PS=1.325 NRD=2.9353 NRS=1.9503 M=1
+ R=6.66667 SA=75001.1 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1003 N_GCLK_M1003_d N_A_1041_387#_M1003_g N_VPWR_M1009_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.530045 PD=1.42 PS=2.2083 NRD=1.7533 NRS=7.0329 M=1
+ R=7.46667 SA=75002 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1005 N_GCLK_M1003_d N_A_1041_387#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=14.4324 P=20.08
*
.include "sky130_fd_sc_hs__dlclkp_2.pxi.spice"
*
.ends
*
*
