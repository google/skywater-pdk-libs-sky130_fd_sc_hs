* File: sky130_fd_sc_hs__a21o_1.pxi.spice
* Created: Tue Sep  1 19:49:34 2020
* 
x_PM_SKY130_FD_SC_HS__A21O_1%A_81_264# N_A_81_264#_M1006_d N_A_81_264#_M1001_s
+ N_A_81_264#_c_60_n N_A_81_264#_M1000_g N_A_81_264#_c_61_n N_A_81_264#_c_62_n
+ N_A_81_264#_M1004_g N_A_81_264#_c_63_n N_A_81_264#_c_67_n N_A_81_264#_c_71_p
+ N_A_81_264#_c_64_n N_A_81_264#_c_65_n N_A_81_264#_c_68_n N_A_81_264#_c_69_n
+ PM_SKY130_FD_SC_HS__A21O_1%A_81_264#
x_PM_SKY130_FD_SC_HS__A21O_1%B1 N_B1_c_121_n N_B1_M1001_g N_B1_M1006_g B1
+ PM_SKY130_FD_SC_HS__A21O_1%B1
x_PM_SKY130_FD_SC_HS__A21O_1%A1 N_A1_M1007_g N_A1_c_153_n N_A1_M1003_g A1
+ PM_SKY130_FD_SC_HS__A21O_1%A1
x_PM_SKY130_FD_SC_HS__A21O_1%A2 N_A2_M1005_g N_A2_c_187_n N_A2_c_188_n
+ N_A2_c_193_n N_A2_M1002_g N_A2_c_189_n A2 N_A2_c_191_n
+ PM_SKY130_FD_SC_HS__A21O_1%A2
x_PM_SKY130_FD_SC_HS__A21O_1%X N_X_M1004_s N_X_M1000_s N_X_c_222_n N_X_c_223_n
+ N_X_c_224_n X X X X N_X_c_225_n PM_SKY130_FD_SC_HS__A21O_1%X
x_PM_SKY130_FD_SC_HS__A21O_1%VPWR N_VPWR_M1000_d N_VPWR_M1003_d N_VPWR_c_243_n
+ N_VPWR_c_244_n N_VPWR_c_245_n N_VPWR_c_246_n VPWR N_VPWR_c_247_n
+ N_VPWR_c_248_n N_VPWR_c_242_n N_VPWR_c_250_n PM_SKY130_FD_SC_HS__A21O_1%VPWR
x_PM_SKY130_FD_SC_HS__A21O_1%A_364_392# N_A_364_392#_M1001_d
+ N_A_364_392#_M1002_d N_A_364_392#_c_278_n N_A_364_392#_c_279_n
+ N_A_364_392#_c_280_n N_A_364_392#_c_281_n N_A_364_392#_c_282_n
+ PM_SKY130_FD_SC_HS__A21O_1%A_364_392#
x_PM_SKY130_FD_SC_HS__A21O_1%VGND N_VGND_M1004_d N_VGND_M1005_d N_VGND_c_309_n
+ N_VGND_c_310_n N_VGND_c_343_n N_VGND_c_335_n N_VGND_c_311_n N_VGND_c_312_n
+ N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n VGND N_VGND_c_316_n
+ N_VGND_c_317_n PM_SKY130_FD_SC_HS__A21O_1%VGND
cc_1 VNB N_A_81_264#_c_60_n 0.0396791f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_2 VNB N_A_81_264#_c_61_n 0.03594f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.47
cc_3 VNB N_A_81_264#_c_62_n 0.0196825f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.395
cc_4 VNB N_A_81_264#_c_63_n 0.0196318f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.485
cc_5 VNB N_A_81_264#_c_64_n 0.00381609f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=0.805
cc_6 VNB N_A_81_264#_c_65_n 0.00278456f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.38
cc_7 VNB N_B1_c_121_n 0.0197428f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=0.68
cc_8 VNB N_B1_M1006_g 0.0197271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB B1 8.71858e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_10 VNB N_A1_M1007_g 0.0191344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_153_n 0.0194427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A1 0.0032213f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_13 VNB N_A2_M1005_g 0.012615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_187_n 0.00849485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_188_n 0.0145107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_189_n 0.050643f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.95
cc_17 VNB A2 0.0277287f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_18 VNB N_A2_c_191_n 5.28587e-19 $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.815
cc_19 VNB N_X_c_222_n 0.0282147f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_20 VNB N_X_c_223_n 0.0149129f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.47
cc_21 VNB N_X_c_224_n 0.0121113f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.95
cc_22 VNB N_X_c_225_n 0.0283359f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.115
cc_23 VNB N_VPWR_c_242_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.47
cc_24 VNB N_VGND_c_309_n 0.0280514f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_25 VNB N_VGND_c_310_n 0.0219582f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.395
cc_26 VNB N_VGND_c_311_n 0.0410501f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_27 VNB N_VGND_c_312_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_28 VNB N_VGND_c_313_n 0.0214589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_314_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.65
cc_30 VNB N_VGND_c_315_n 0.0245056f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.95
cc_31 VNB N_VGND_c_316_n 0.0245652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_317_n 0.243932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A_81_264#_c_60_n 0.0295754f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_34 VPB N_A_81_264#_c_67_n 0.0167758f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.815
cc_35 VPB N_A_81_264#_c_68_n 0.00511476f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.115
cc_36 VPB N_A_81_264#_c_69_n 0.00741545f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.95
cc_37 VPB N_B1_c_121_n 0.0399964f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.68
cc_38 VPB B1 0.00206873f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_39 VPB N_A1_c_153_n 0.0355337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB A1 0.00137164f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_41 VPB N_A2_c_188_n 0.0112268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A2_c_193_n 0.0297875f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_43 VPB X 0.00942864f $X=-0.19 $Y=1.66 $X2=1.245 $Y2=1.485
cc_44 VPB X 0.0420202f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.815
cc_45 VPB N_X_c_225_n 0.00787925f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=2.115
cc_46 VPB N_VPWR_c_243_n 0.029481f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_47 VPB N_VPWR_c_244_n 0.00835244f $X=-0.19 $Y=1.66 $X2=1.245 $Y2=1.485
cc_48 VPB N_VPWR_c_245_n 0.0407193f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_49 VPB N_VPWR_c_246_n 0.00382106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_247_n 0.0196317f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=2.13
cc_51 VPB N_VPWR_c_248_n 0.0258341f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.95
cc_52 VPB N_VPWR_c_242_n 0.0875264f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.47
cc_53 VPB N_VPWR_c_250_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_364_392#_c_278_n 0.00419085f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_55 VPB N_A_364_392#_c_279_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_56 VPB N_A_364_392#_c_280_n 0.00800581f $X=-0.19 $Y=1.66 $X2=0.755 $Y2=1.47
cc_57 VPB N_A_364_392#_c_281_n 0.0133173f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.95
cc_58 VPB N_A_364_392#_c_282_n 0.0360166f $X=-0.19 $Y=1.66 $X2=1.245 $Y2=1.485
cc_59 N_A_81_264#_c_61_n N_B1_c_121_n 0.00540357f $X=1.13 $Y=1.47 $X2=-0.19
+ $Y2=-0.245
cc_60 N_A_81_264#_c_71_p N_B1_c_121_n 0.00275112f $X=1.805 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_61 N_A_81_264#_c_65_n N_B1_c_121_n 0.00340356f $X=1.33 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_62 N_A_81_264#_c_68_n N_B1_c_121_n 0.00700954f $X=1.52 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_63 N_A_81_264#_c_69_n N_B1_c_121_n 0.00860612f $X=1.425 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_64 N_A_81_264#_c_62_n N_B1_M1006_g 0.0176258f $X=1.205 $Y=1.395 $X2=0 $Y2=0
cc_65 N_A_81_264#_c_71_p N_B1_M1006_g 0.0121724f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_66 N_A_81_264#_c_64_n N_B1_M1006_g 0.00723827f $X=1.97 $Y=0.805 $X2=0 $Y2=0
cc_67 N_A_81_264#_c_65_n N_B1_M1006_g 0.00411569f $X=1.33 $Y=1.38 $X2=0 $Y2=0
cc_68 N_A_81_264#_c_71_p B1 0.0159378f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_69 N_A_81_264#_c_65_n B1 0.0165507f $X=1.33 $Y=1.38 $X2=0 $Y2=0
cc_70 N_A_81_264#_c_68_n B1 0.00152541f $X=1.52 $Y=2.115 $X2=0 $Y2=0
cc_71 N_A_81_264#_c_69_n B1 0.00952856f $X=1.425 $Y=1.95 $X2=0 $Y2=0
cc_72 N_A_81_264#_c_71_p N_A1_M1007_g 0.00346932f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_73 N_A_81_264#_c_64_n N_A1_M1007_g 0.00599966f $X=1.97 $Y=0.805 $X2=0 $Y2=0
cc_74 N_A_81_264#_c_71_p N_A1_c_153_n 3.32928e-19 $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_75 N_A_81_264#_c_71_p A1 0.00468798f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_76 N_A_81_264#_c_71_p N_A2_M1005_g 5.14251e-19 $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_77 N_A_81_264#_c_64_n N_A2_M1005_g 4.72693e-19 $X=1.97 $Y=0.805 $X2=0 $Y2=0
cc_78 N_A_81_264#_c_60_n N_X_c_222_n 0.00857934f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_81_264#_c_61_n N_X_c_222_n 0.00199362f $X=1.13 $Y=1.47 $X2=0 $Y2=0
cc_80 N_A_81_264#_c_63_n N_X_c_222_n 0.0514037f $X=1.245 $Y=1.485 $X2=0 $Y2=0
cc_81 N_A_81_264#_c_60_n X 0.00308687f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_81_264#_c_63_n X 7.18422e-19 $X=1.245 $Y=1.485 $X2=0 $Y2=0
cc_83 N_A_81_264#_c_60_n X 0.0121388f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_81_264#_c_60_n N_X_c_225_n 0.0142219f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_81_264#_c_63_n N_X_c_225_n 0.0262118f $X=1.245 $Y=1.485 $X2=0 $Y2=0
cc_86 N_A_81_264#_c_60_n N_VPWR_c_243_n 0.0128637f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_81_264#_c_61_n N_VPWR_c_243_n 7.91918e-19 $X=1.13 $Y=1.47 $X2=0 $Y2=0
cc_88 N_A_81_264#_c_63_n N_VPWR_c_243_n 0.0214461f $X=1.245 $Y=1.485 $X2=0 $Y2=0
cc_89 N_A_81_264#_c_69_n N_VPWR_c_243_n 0.0563013f $X=1.425 $Y=1.95 $X2=0 $Y2=0
cc_90 N_A_81_264#_c_67_n N_VPWR_c_245_n 0.0159743f $X=1.52 $Y=2.815 $X2=0 $Y2=0
cc_91 N_A_81_264#_c_60_n N_VPWR_c_247_n 0.00445602f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_92 N_A_81_264#_c_60_n N_VPWR_c_242_n 0.00865852f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_93 N_A_81_264#_c_67_n N_VPWR_c_242_n 0.0132221f $X=1.52 $Y=2.815 $X2=0 $Y2=0
cc_94 N_A_81_264#_c_71_p N_A_364_392#_c_278_n 0.00628732f $X=1.805 $Y=1.195
+ $X2=0 $Y2=0
cc_95 N_A_81_264#_c_68_n N_A_364_392#_c_278_n 0.0124439f $X=1.52 $Y=2.115 $X2=0
+ $Y2=0
cc_96 N_A_81_264#_c_68_n N_A_364_392#_c_279_n 0.059268f $X=1.52 $Y=2.115 $X2=0
+ $Y2=0
cc_97 N_A_81_264#_c_71_p N_VGND_M1004_d 0.00682387f $X=1.805 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_81_264#_c_65_n N_VGND_M1004_d 0.00136247f $X=1.33 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_81_264#_c_62_n N_VGND_c_309_n 0.0157678f $X=1.205 $Y=1.395 $X2=0 $Y2=0
cc_100 N_A_81_264#_c_71_p N_VGND_c_309_n 0.0137131f $X=1.805 $Y=1.195 $X2=0
+ $Y2=0
cc_101 N_A_81_264#_c_64_n N_VGND_c_309_n 0.0178602f $X=1.97 $Y=0.805 $X2=0 $Y2=0
cc_102 N_A_81_264#_c_65_n N_VGND_c_309_n 0.00902191f $X=1.33 $Y=1.38 $X2=0 $Y2=0
cc_103 N_A_81_264#_c_64_n N_VGND_c_310_n 0.00746887f $X=1.97 $Y=0.805 $X2=0
+ $Y2=0
cc_104 N_A_81_264#_c_62_n N_VGND_c_311_n 0.00365567f $X=1.205 $Y=1.395 $X2=0
+ $Y2=0
cc_105 N_A_81_264#_c_64_n N_VGND_c_313_n 0.00615803f $X=1.97 $Y=0.805 $X2=0
+ $Y2=0
cc_106 N_A_81_264#_c_71_p N_VGND_c_315_n 0.00495397f $X=1.805 $Y=1.195 $X2=0
+ $Y2=0
cc_107 N_A_81_264#_c_64_n N_VGND_c_315_n 0.00276199f $X=1.97 $Y=0.805 $X2=0
+ $Y2=0
cc_108 N_A_81_264#_c_62_n N_VGND_c_317_n 0.00404919f $X=1.205 $Y=1.395 $X2=0
+ $Y2=0
cc_109 N_A_81_264#_c_64_n N_VGND_c_317_n 0.00967008f $X=1.97 $Y=0.805 $X2=0
+ $Y2=0
cc_110 N_B1_M1006_g N_A1_M1007_g 0.0117284f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_111 N_B1_c_121_n N_A1_c_153_n 0.0345548f $X=1.745 $Y=1.885 $X2=0 $Y2=0
cc_112 B1 N_A1_c_153_n 0.00115083f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_113 N_B1_c_121_n A1 0.00114936f $X=1.745 $Y=1.885 $X2=0 $Y2=0
cc_114 B1 A1 0.0204777f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_115 N_B1_c_121_n N_VPWR_c_245_n 0.00445602f $X=1.745 $Y=1.885 $X2=0 $Y2=0
cc_116 N_B1_c_121_n N_VPWR_c_242_n 0.00863237f $X=1.745 $Y=1.885 $X2=0 $Y2=0
cc_117 N_B1_c_121_n N_A_364_392#_c_278_n 0.00261932f $X=1.745 $Y=1.885 $X2=0
+ $Y2=0
cc_118 B1 N_A_364_392#_c_278_n 0.00238988f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_119 N_B1_c_121_n N_A_364_392#_c_279_n 0.00960248f $X=1.745 $Y=1.885 $X2=0
+ $Y2=0
cc_120 N_B1_M1006_g N_VGND_c_309_n 0.00552238f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_121 N_B1_M1006_g N_VGND_c_313_n 0.0037378f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_122 N_B1_M1006_g N_VGND_c_317_n 0.00454494f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_123 N_A1_c_153_n N_A2_c_187_n 0.0214073f $X=2.195 $Y=1.885 $X2=0 $Y2=0
cc_124 A1 N_A2_c_187_n 0.00223091f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A1_c_153_n N_A2_c_188_n 0.00512744f $X=2.195 $Y=1.885 $X2=0 $Y2=0
cc_126 N_A1_c_153_n N_A2_c_193_n 0.0172837f $X=2.195 $Y=1.885 $X2=0 $Y2=0
cc_127 N_A1_M1007_g N_A2_c_189_n 0.0301488f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_128 N_A1_c_153_n N_VPWR_c_244_n 0.00507786f $X=2.195 $Y=1.885 $X2=0 $Y2=0
cc_129 N_A1_c_153_n N_VPWR_c_245_n 0.00445602f $X=2.195 $Y=1.885 $X2=0 $Y2=0
cc_130 N_A1_c_153_n N_VPWR_c_242_n 0.0085802f $X=2.195 $Y=1.885 $X2=0 $Y2=0
cc_131 N_A1_c_153_n N_A_364_392#_c_278_n 0.00146854f $X=2.195 $Y=1.885 $X2=0
+ $Y2=0
cc_132 A1 N_A_364_392#_c_278_n 0.00747456f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A1_c_153_n N_A_364_392#_c_279_n 0.0104821f $X=2.195 $Y=1.885 $X2=0
+ $Y2=0
cc_134 N_A1_c_153_n N_A_364_392#_c_280_n 0.0131434f $X=2.195 $Y=1.885 $X2=0
+ $Y2=0
cc_135 A1 N_A_364_392#_c_280_n 0.0175118f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A1_c_153_n N_A_364_392#_c_282_n 6.36743e-19 $X=2.195 $Y=1.885 $X2=0
+ $Y2=0
cc_137 N_A1_M1007_g N_VGND_c_310_n 0.00365891f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_138 N_A1_c_153_n N_VGND_c_335_n 4.2417e-19 $X=2.195 $Y=1.885 $X2=0 $Y2=0
cc_139 A1 N_VGND_c_335_n 0.00247219f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_140 N_A1_M1007_g N_VGND_c_313_n 0.0037378f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_141 N_A1_M1007_g N_VGND_c_315_n 0.00110784f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_142 N_A1_M1007_g N_VGND_c_317_n 0.00454494f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_143 N_A2_c_193_n N_VPWR_c_244_n 0.00507786f $X=2.675 $Y=1.885 $X2=0 $Y2=0
cc_144 N_A2_c_193_n N_VPWR_c_248_n 0.00445602f $X=2.675 $Y=1.885 $X2=0 $Y2=0
cc_145 N_A2_c_193_n N_VPWR_c_242_n 0.00861892f $X=2.675 $Y=1.885 $X2=0 $Y2=0
cc_146 N_A2_c_193_n N_A_364_392#_c_279_n 6.36743e-19 $X=2.675 $Y=1.885 $X2=0
+ $Y2=0
cc_147 N_A2_c_193_n N_A_364_392#_c_280_n 0.0165246f $X=2.675 $Y=1.885 $X2=0
+ $Y2=0
cc_148 N_A2_c_193_n N_A_364_392#_c_281_n 0.0017173f $X=2.675 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_A2_c_193_n N_A_364_392#_c_282_n 0.0106338f $X=2.675 $Y=1.885 $X2=0
+ $Y2=0
cc_150 N_A2_c_189_n N_VGND_c_310_n 0.0130563f $X=2.81 $Y=0.405 $X2=0 $Y2=0
cc_151 A2 N_VGND_c_310_n 0.0034499f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_152 N_A2_c_191_n N_VGND_c_310_n 0.02473f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_153 N_A2_M1005_g N_VGND_c_343_n 0.0124199f $X=2.66 $Y=1 $X2=0 $Y2=0
cc_154 N_A2_c_191_n N_VGND_c_343_n 0.0029673f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_155 N_A2_M1005_g N_VGND_c_315_n 0.0103623f $X=2.66 $Y=1 $X2=0 $Y2=0
cc_156 N_A2_c_187_n N_VGND_c_315_n 0.00110067f $X=2.675 $Y=1.485 $X2=0 $Y2=0
cc_157 N_A2_c_189_n N_VGND_c_315_n 0.0050123f $X=2.81 $Y=0.405 $X2=0 $Y2=0
cc_158 A2 N_VGND_c_315_n 0.00291185f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_159 N_A2_c_191_n N_VGND_c_315_n 0.0137799f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_160 N_A2_c_189_n N_VGND_c_316_n 0.00760015f $X=2.81 $Y=0.405 $X2=0 $Y2=0
cc_161 N_A2_c_191_n N_VGND_c_316_n 0.0389306f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_162 N_A2_c_189_n N_VGND_c_317_n 0.00934546f $X=2.81 $Y=0.405 $X2=0 $Y2=0
cc_163 N_A2_c_191_n N_VGND_c_317_n 0.0210356f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_164 X N_VPWR_c_243_n 0.0781509f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_165 X N_VPWR_c_247_n 0.0154862f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_166 X N_VPWR_c_242_n 0.0127853f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_167 N_X_c_224_n N_VGND_c_311_n 0.00435429f $X=0.99 $Y=0.885 $X2=0 $Y2=0
cc_168 N_X_c_224_n N_VGND_c_317_n 0.00720812f $X=0.99 $Y=0.885 $X2=0 $Y2=0
cc_169 N_VPWR_c_244_n N_A_364_392#_c_279_n 0.0455206f $X=2.435 $Y=2.455 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_245_n N_A_364_392#_c_279_n 0.014552f $X=2.335 $Y=3.33 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_242_n N_A_364_392#_c_279_n 0.0119791f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_172 N_VPWR_M1003_d N_A_364_392#_c_280_n 0.00279158f $X=2.27 $Y=1.96 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_244_n N_A_364_392#_c_280_n 0.016109f $X=2.435 $Y=2.455 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_244_n N_A_364_392#_c_282_n 0.0455206f $X=2.435 $Y=2.455 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_248_n N_A_364_392#_c_282_n 0.0145938f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_242_n N_A_364_392#_c_282_n 0.0120466f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_177 N_A_364_392#_c_280_n N_VGND_c_315_n 6.04679e-19 $X=2.735 $Y=2.035 $X2=0
+ $Y2=0
cc_178 N_A_364_392#_c_281_n N_VGND_c_315_n 0.0114345f $X=2.9 $Y=2.12 $X2=0 $Y2=0
cc_179 N_VGND_c_310_n A_452_136# 0.00255642f $X=2.39 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_180 N_VGND_c_343_n A_452_136# 0.00302954f $X=2.71 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_181 N_VGND_c_335_n A_452_136# 0.00617481f $X=2.475 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
