* File: sky130_fd_sc_hs__sdfrtp_4.pxi.spice
* Created: Thu Aug 27 21:08:59 2020
* 
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_27_74# N_A_27_74#_M1037_s N_A_27_74#_M1021_s
+ N_A_27_74#_c_299_n N_A_27_74#_c_300_n N_A_27_74#_M1009_g N_A_27_74#_c_306_n
+ N_A_27_74#_M1036_g N_A_27_74#_c_301_n N_A_27_74#_c_302_n N_A_27_74#_c_308_n
+ N_A_27_74#_c_303_n N_A_27_74#_c_309_n N_A_27_74#_c_304_n N_A_27_74#_c_310_n
+ N_A_27_74#_c_311_n N_A_27_74#_c_305_n PM_SKY130_FD_SC_HS__SDFRTP_4%A_27_74#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%SCE N_SCE_c_390_n N_SCE_M1037_g N_SCE_c_391_n
+ N_SCE_M1021_g N_SCE_c_392_n N_SCE_c_393_n N_SCE_M1017_g N_SCE_c_382_n
+ N_SCE_M1039_g N_SCE_c_384_n N_SCE_c_385_n N_SCE_c_386_n N_SCE_c_387_n SCE SCE
+ SCE N_SCE_c_388_n SCE N_SCE_c_389_n PM_SKY130_FD_SC_HS__SDFRTP_4%SCE
x_PM_SKY130_FD_SC_HS__SDFRTP_4%D N_D_M1010_g N_D_c_470_n N_D_c_475_n N_D_M1033_g
+ D N_D_c_471_n N_D_c_472_n N_D_c_473_n PM_SKY130_FD_SC_HS__SDFRTP_4%D
x_PM_SKY130_FD_SC_HS__SDFRTP_4%SCD N_SCD_c_520_n N_SCD_M1006_g N_SCD_M1040_g
+ N_SCD_c_517_n SCD SCD N_SCD_c_519_n PM_SKY130_FD_SC_HS__SDFRTP_4%SCD
x_PM_SKY130_FD_SC_HS__SDFRTP_4%RESET_B N_RESET_B_M1023_g N_RESET_B_c_569_n
+ N_RESET_B_M1045_g N_RESET_B_c_563_n N_RESET_B_M1030_g N_RESET_B_c_564_n
+ N_RESET_B_c_565_n N_RESET_B_c_570_n N_RESET_B_M1020_g N_RESET_B_c_566_n
+ N_RESET_B_M1041_g N_RESET_B_c_573_n N_RESET_B_c_574_n N_RESET_B_M1038_g
+ N_RESET_B_c_575_n N_RESET_B_c_576_n N_RESET_B_c_577_n N_RESET_B_c_578_n
+ N_RESET_B_c_579_n RESET_B N_RESET_B_c_581_n N_RESET_B_c_582_n
+ N_RESET_B_c_583_n N_RESET_B_c_584_n N_RESET_B_c_585_n
+ PM_SKY130_FD_SC_HS__SDFRTP_4%RESET_B
x_PM_SKY130_FD_SC_HS__SDFRTP_4%CLK N_CLK_c_768_n N_CLK_M1019_g N_CLK_M1007_g
+ N_CLK_c_770_n N_CLK_c_781_n CLK N_CLK_c_771_n PM_SKY130_FD_SC_HS__SDFRTP_4%CLK
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_1034_74# N_A_1034_74#_M1015_d
+ N_A_1034_74#_M1031_d N_A_1034_74#_c_844_n N_A_1034_74#_c_845_n
+ N_A_1034_74#_M1046_g N_A_1034_74#_c_823_n N_A_1034_74#_M1016_g
+ N_A_1034_74#_c_825_n N_A_1034_74#_M1008_g N_A_1034_74#_c_826_n
+ N_A_1034_74#_c_827_n N_A_1034_74#_c_847_n N_A_1034_74#_M1043_g
+ N_A_1034_74#_c_828_n N_A_1034_74#_c_829_n N_A_1034_74#_c_830_n
+ N_A_1034_74#_c_831_n N_A_1034_74#_c_832_n N_A_1034_74#_c_833_n
+ N_A_1034_74#_c_858_n N_A_1034_74#_c_834_n N_A_1034_74#_c_835_n
+ N_A_1034_74#_c_836_n N_A_1034_74#_c_837_n N_A_1034_74#_c_860_n
+ N_A_1034_74#_c_850_n N_A_1034_74#_c_838_n N_A_1034_74#_c_839_n
+ N_A_1034_74#_c_840_n N_A_1034_74#_c_841_n N_A_1034_74#_c_842_n
+ N_A_1034_74#_c_843_n PM_SKY130_FD_SC_HS__SDFRTP_4%A_1034_74#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_1367_112# N_A_1367_112#_M1025_d
+ N_A_1367_112#_M1000_d N_A_1367_112#_M1001_g N_A_1367_112#_c_1048_n
+ N_A_1367_112#_c_1049_n N_A_1367_112#_M1032_g N_A_1367_112#_c_1044_n
+ N_A_1367_112#_c_1045_n N_A_1367_112#_c_1067_n N_A_1367_112#_c_1046_n
+ N_A_1367_112#_c_1047_n N_A_1367_112#_c_1053_n N_A_1367_112#_c_1070_n
+ N_A_1367_112#_c_1094_n PM_SKY130_FD_SC_HS__SDFRTP_4%A_1367_112#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_1233_138# N_A_1233_138#_M1024_d
+ N_A_1233_138#_M1046_d N_A_1233_138#_M1020_d N_A_1233_138#_M1025_g
+ N_A_1233_138#_c_1153_n N_A_1233_138#_c_1161_n N_A_1233_138#_M1000_g
+ N_A_1233_138#_c_1162_n N_A_1233_138#_c_1171_n N_A_1233_138#_c_1154_n
+ N_A_1233_138#_c_1174_n N_A_1233_138#_c_1155_n N_A_1233_138#_c_1156_n
+ N_A_1233_138#_c_1157_n N_A_1233_138#_c_1158_n N_A_1233_138#_c_1159_n
+ N_A_1233_138#_c_1166_n PM_SKY130_FD_SC_HS__SDFRTP_4%A_1233_138#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_855_368# N_A_855_368#_M1007_s
+ N_A_855_368#_M1019_s N_A_855_368#_c_1287_n N_A_855_368#_M1015_g
+ N_A_855_368#_c_1288_n N_A_855_368#_M1031_g N_A_855_368#_c_1289_n
+ N_A_855_368#_c_1290_n N_A_855_368#_c_1291_n N_A_855_368#_c_1303_n
+ N_A_855_368#_c_1304_n N_A_855_368#_c_1292_n N_A_855_368#_M1024_g
+ N_A_855_368#_c_1305_n N_A_855_368#_c_1306_n N_A_855_368#_c_1307_n
+ N_A_855_368#_M1042_g N_A_855_368#_c_1308_n N_A_855_368#_c_1309_n
+ N_A_855_368#_c_1310_n N_A_855_368#_M1003_g N_A_855_368#_c_1293_n
+ N_A_855_368#_c_1294_n N_A_855_368#_M1034_g N_A_855_368#_c_1296_n
+ N_A_855_368#_c_1314_n N_A_855_368#_c_1297_n N_A_855_368#_c_1339_n
+ N_A_855_368#_c_1326_n N_A_855_368#_c_1315_n N_A_855_368#_c_1298_n
+ N_A_855_368#_c_1299_n N_A_855_368#_c_1317_n N_A_855_368#_c_1300_n
+ PM_SKY130_FD_SC_HS__SDFRTP_4%A_855_368#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_2003_48# N_A_2003_48#_M1027_d
+ N_A_2003_48#_M1038_d N_A_2003_48#_M1028_g N_A_2003_48#_c_1485_n
+ N_A_2003_48#_c_1494_n N_A_2003_48#_M1026_g N_A_2003_48#_c_1486_n
+ N_A_2003_48#_c_1487_n N_A_2003_48#_c_1488_n N_A_2003_48#_c_1489_n
+ N_A_2003_48#_c_1490_n N_A_2003_48#_c_1495_n N_A_2003_48#_c_1491_n
+ N_A_2003_48#_c_1492_n PM_SKY130_FD_SC_HS__SDFRTP_4%A_2003_48#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_1745_74# N_A_1745_74#_M1008_d
+ N_A_1745_74#_M1003_d N_A_1745_74#_c_1573_n N_A_1745_74#_M1027_g
+ N_A_1745_74#_c_1574_n N_A_1745_74#_c_1589_n N_A_1745_74#_c_1590_n
+ N_A_1745_74#_M1022_g N_A_1745_74#_c_1575_n N_A_1745_74#_c_1591_n
+ N_A_1745_74#_M1012_g N_A_1745_74#_c_1576_n N_A_1745_74#_M1013_g
+ N_A_1745_74#_c_1577_n N_A_1745_74#_c_1578_n N_A_1745_74#_c_1593_n
+ N_A_1745_74#_M1014_g N_A_1745_74#_c_1579_n N_A_1745_74#_c_1580_n
+ N_A_1745_74#_c_1581_n N_A_1745_74#_c_1626_n N_A_1745_74#_c_1595_n
+ N_A_1745_74#_c_1582_n N_A_1745_74#_c_1583_n N_A_1745_74#_c_1584_n
+ N_A_1745_74#_c_1597_n N_A_1745_74#_c_1598_n N_A_1745_74#_c_1599_n
+ N_A_1745_74#_c_1585_n N_A_1745_74#_c_1586_n N_A_1745_74#_c_1587_n
+ PM_SKY130_FD_SC_HS__SDFRTP_4%A_1745_74#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_2339_74# N_A_2339_74#_M1013_s
+ N_A_2339_74#_M1012_d N_A_2339_74#_c_1737_n N_A_2339_74#_M1011_g
+ N_A_2339_74#_c_1738_n N_A_2339_74#_c_1739_n N_A_2339_74#_c_1740_n
+ N_A_2339_74#_M1018_g N_A_2339_74#_c_1748_n N_A_2339_74#_M1002_g
+ N_A_2339_74#_c_1749_n N_A_2339_74#_M1004_g N_A_2339_74#_c_1750_n
+ N_A_2339_74#_M1005_g N_A_2339_74#_c_1741_n N_A_2339_74#_M1029_g
+ N_A_2339_74#_c_1751_n N_A_2339_74#_M1044_g N_A_2339_74#_c_1742_n
+ N_A_2339_74#_M1035_g N_A_2339_74#_c_1743_n N_A_2339_74#_c_1744_n
+ N_A_2339_74#_c_1745_n N_A_2339_74#_c_1746_n N_A_2339_74#_c_1747_n
+ PM_SKY130_FD_SC_HS__SDFRTP_4%A_2339_74#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%VPWR N_VPWR_M1021_d N_VPWR_M1006_d N_VPWR_M1019_d
+ N_VPWR_M1032_d N_VPWR_M1000_s N_VPWR_M1026_d N_VPWR_M1022_d N_VPWR_M1014_s
+ N_VPWR_M1004_d N_VPWR_M1044_d N_VPWR_c_1855_n N_VPWR_c_1856_n N_VPWR_c_1857_n
+ N_VPWR_c_1858_n N_VPWR_c_1859_n N_VPWR_c_1860_n N_VPWR_c_1861_n
+ N_VPWR_c_1862_n N_VPWR_c_1863_n N_VPWR_c_1864_n N_VPWR_c_1865_n
+ N_VPWR_c_1866_n N_VPWR_c_1867_n N_VPWR_c_1868_n N_VPWR_c_1869_n
+ N_VPWR_c_1870_n VPWR N_VPWR_c_1871_n N_VPWR_c_1872_n N_VPWR_c_1873_n
+ N_VPWR_c_1874_n N_VPWR_c_1875_n N_VPWR_c_1876_n N_VPWR_c_1877_n
+ N_VPWR_c_1878_n N_VPWR_c_1879_n N_VPWR_c_1880_n N_VPWR_c_1881_n
+ N_VPWR_c_1882_n N_VPWR_c_1883_n N_VPWR_c_1854_n
+ PM_SKY130_FD_SC_HS__SDFRTP_4%VPWR
x_PM_SKY130_FD_SC_HS__SDFRTP_4%A_415_81# N_A_415_81#_M1010_d N_A_415_81#_M1024_s
+ N_A_415_81#_M1033_d N_A_415_81#_M1045_d N_A_415_81#_M1046_s
+ N_A_415_81#_c_2044_n N_A_415_81#_c_2059_n N_A_415_81#_c_2045_n
+ N_A_415_81#_c_2046_n N_A_415_81#_c_2052_n N_A_415_81#_c_2053_n
+ N_A_415_81#_c_2054_n N_A_415_81#_c_2047_n N_A_415_81#_c_2048_n
+ N_A_415_81#_c_2049_n N_A_415_81#_c_2055_n N_A_415_81#_c_2050_n
+ N_A_415_81#_c_2057_n N_A_415_81#_c_2058_n
+ PM_SKY130_FD_SC_HS__SDFRTP_4%A_415_81#
x_PM_SKY130_FD_SC_HS__SDFRTP_4%Q N_Q_M1011_s N_Q_M1029_s N_Q_M1002_s N_Q_M1005_s
+ N_Q_c_2193_n N_Q_c_2204_n N_Q_c_2208_n N_Q_c_2197_n N_Q_c_2198_n N_Q_c_2199_n
+ N_Q_c_2200_n N_Q_c_2194_n N_Q_c_2195_n Q PM_SKY130_FD_SC_HS__SDFRTP_4%Q
x_PM_SKY130_FD_SC_HS__SDFRTP_4%VGND N_VGND_M1037_d N_VGND_M1023_d N_VGND_M1007_d
+ N_VGND_M1030_d N_VGND_M1028_d N_VGND_M1013_d N_VGND_M1018_d N_VGND_M1035_d
+ N_VGND_c_2260_n N_VGND_c_2261_n N_VGND_c_2262_n N_VGND_c_2263_n
+ N_VGND_c_2264_n N_VGND_c_2265_n N_VGND_c_2266_n N_VGND_c_2267_n
+ N_VGND_c_2268_n N_VGND_c_2269_n N_VGND_c_2270_n VGND N_VGND_c_2271_n
+ N_VGND_c_2272_n N_VGND_c_2273_n N_VGND_c_2274_n N_VGND_c_2275_n
+ N_VGND_c_2276_n N_VGND_c_2277_n N_VGND_c_2278_n N_VGND_c_2279_n
+ N_VGND_c_2280_n N_VGND_c_2281_n N_VGND_c_2282_n
+ PM_SKY130_FD_SC_HS__SDFRTP_4%VGND
x_PM_SKY130_FD_SC_HS__SDFRTP_4%noxref_24 N_noxref_24_M1009_s N_noxref_24_M1040_d
+ N_noxref_24_c_2403_n N_noxref_24_c_2404_n N_noxref_24_c_2405_n
+ PM_SKY130_FD_SC_HS__SDFRTP_4%noxref_24
cc_1 VNB N_A_27_74#_c_299_n 0.0258189f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_2 VNB N_A_27_74#_c_300_n 0.0213547f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_3 VNB N_A_27_74#_c_301_n 0.0257773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_4 VNB N_A_27_74#_c_302_n 0.0190417f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_5 VNB N_A_27_74#_c_303_n 0.00987534f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_6 VNB N_A_27_74#_c_304_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_7 VNB N_A_27_74#_c_305_n 0.0395906f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_8 VNB N_SCE_M1037_g 0.0668709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_c_382_n 0.0578303f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_10 VNB N_SCE_M1039_g 0.0224937f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_11 VNB N_SCE_c_384_n 0.00775502f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_12 VNB N_SCE_c_385_n 0.0420954f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_13 VNB N_SCE_c_386_n 0.0131161f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_14 VNB N_SCE_c_387_n 0.00292005f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_15 VNB N_SCE_c_388_n 0.0106235f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_16 VNB N_SCE_c_389_n 0.00168276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_c_470_n 0.0279786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_D_c_471_n 0.0381417f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.245
cc_19 VNB N_D_c_472_n 0.00727955f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_20 VNB N_D_c_473_n 0.0173744f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_21 VNB N_SCD_M1040_g 0.0408649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCD_c_517_n 0.00419656f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_23 VNB SCD 0.00223563f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_24 VNB N_SCD_c_519_n 0.0167355f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_25 VNB N_RESET_B_M1023_g 0.0595346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_RESET_B_c_563_n 0.0177368f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.01
cc_27 VNB N_RESET_B_c_564_n 0.0238599f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_28 VNB N_RESET_B_c_565_n 0.00691999f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.245
cc_29 VNB N_RESET_B_c_566_n 0.0181108f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_30 VNB N_RESET_B_M1041_g 0.0569134f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_31 VNB N_CLK_c_768_n 0.0191031f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_32 VNB N_CLK_M1007_g 0.022731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_CLK_c_770_n 0.0606573f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_34 VNB N_CLK_c_771_n 0.0108773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_35 VNB N_A_1034_74#_c_823_n 0.00940815f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_36 VNB N_A_1034_74#_M1016_g 0.0369745f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_37 VNB N_A_1034_74#_c_825_n 0.0168538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1034_74#_c_826_n 0.0237434f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_39 VNB N_A_1034_74#_c_827_n 0.00657402f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_40 VNB N_A_1034_74#_c_828_n 0.006943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1034_74#_c_829_n 0.00304546f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_42 VNB N_A_1034_74#_c_830_n 0.0383951f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_43 VNB N_A_1034_74#_c_831_n 0.00492357f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_44 VNB N_A_1034_74#_c_832_n 0.00178893f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_45 VNB N_A_1034_74#_c_833_n 0.00102705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1034_74#_c_834_n 0.00657839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1034_74#_c_835_n 0.00231075f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_48 VNB N_A_1034_74#_c_836_n 0.00144678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1034_74#_c_837_n 0.005194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1034_74#_c_838_n 0.00270991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1034_74#_c_839_n 7.04021e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1034_74#_c_840_n 0.0119096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1034_74#_c_841_n 0.0332641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1034_74#_c_842_n 0.00593212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1034_74#_c_843_n 0.00982845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1367_112#_M1001_g 0.0358811f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.935
cc_57 VNB N_A_1367_112#_c_1044_n 0.00473079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1367_112#_c_1045_n 0.0144748f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_59 VNB N_A_1367_112#_c_1046_n 0.00556937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1367_112#_c_1047_n 0.00450848f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.1
cc_61 VNB N_A_1233_138#_M1025_g 0.0225417f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_62 VNB N_A_1233_138#_c_1153_n 0.0164115f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.64
cc_63 VNB N_A_1233_138#_c_1154_n 0.00369363f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_64 VNB N_A_1233_138#_c_1155_n 5.47792e-19 $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_65 VNB N_A_1233_138#_c_1156_n 0.00176601f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.09
cc_66 VNB N_A_1233_138#_c_1157_n 0.00526285f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.09
cc_67 VNB N_A_1233_138#_c_1158_n 0.0281158f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_68 VNB N_A_1233_138#_c_1159_n 0.00236694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_855_368#_c_1287_n 0.0198125f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_70 VNB N_A_855_368#_c_1288_n 0.0327812f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_71 VNB N_A_855_368#_c_1289_n 0.0127252f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_72 VNB N_A_855_368#_c_1290_n 0.0147059f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_73 VNB N_A_855_368#_c_1291_n 0.0254028f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_74 VNB N_A_855_368#_c_1292_n 0.0162132f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_75 VNB N_A_855_368#_c_1293_n 0.019724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_855_368#_c_1294_n 0.00441832f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_77 VNB N_A_855_368#_M1034_g 0.0510568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_855_368#_c_1296_n 0.0072671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_855_368#_c_1297_n 0.00186916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_855_368#_c_1298_n 0.00234418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_855_368#_c_1299_n 0.00183559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_855_368#_c_1300_n 0.00422409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2003_48#_M1028_g 0.0340019f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_84 VNB N_A_2003_48#_c_1485_n 0.0060931f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_85 VNB N_A_2003_48#_c_1486_n 0.0178026f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_86 VNB N_A_2003_48#_c_1487_n 0.00567377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2003_48#_c_1488_n 0.00480935f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_88 VNB N_A_2003_48#_c_1489_n 0.00289977f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_89 VNB N_A_2003_48#_c_1490_n 0.031198f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_90 VNB N_A_2003_48#_c_1491_n 0.00270148f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_91 VNB N_A_2003_48#_c_1492_n 0.00662489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1745_74#_c_1573_n 0.021255f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_93 VNB N_A_1745_74#_c_1574_n 0.00668157f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_94 VNB N_A_1745_74#_c_1575_n 0.0250522f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_95 VNB N_A_1745_74#_c_1576_n 0.0185474f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_96 VNB N_A_1745_74#_c_1577_n 0.0159493f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_97 VNB N_A_1745_74#_c_1578_n 0.014028f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_98 VNB N_A_1745_74#_c_1579_n 0.0143997f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_99 VNB N_A_1745_74#_c_1580_n 0.00251602f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_100 VNB N_A_1745_74#_c_1581_n 0.00496366f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_101 VNB N_A_1745_74#_c_1582_n 0.00146437f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_102 VNB N_A_1745_74#_c_1583_n 0.00359384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1745_74#_c_1584_n 0.0291774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1745_74#_c_1585_n 0.00123798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1745_74#_c_1586_n 0.00179963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1745_74#_c_1587_n 0.0646681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2339_74#_c_1737_n 0.0177259f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_108 VNB N_A_2339_74#_c_1738_n 0.0142247f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_109 VNB N_A_2339_74#_c_1739_n 0.00638412f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_110 VNB N_A_2339_74#_c_1740_n 0.021315f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_111 VNB N_A_2339_74#_c_1741_n 0.0221017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2339_74#_c_1742_n 0.0216728f $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_113 VNB N_A_2339_74#_c_1743_n 0.00311192f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_114 VNB N_A_2339_74#_c_1744_n 0.00104691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2339_74#_c_1745_n 0.00999107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2339_74#_c_1746_n 0.00570341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2339_74#_c_1747_n 0.14135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VPWR_c_1854_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_415_81#_c_2044_n 0.00673461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_415_81#_c_2045_n 0.0163443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_415_81#_c_2046_n 0.00473117f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_122 VNB N_A_415_81#_c_2047_n 0.00322579f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_123 VNB N_A_415_81#_c_2048_n 0.00529525f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_124 VNB N_A_415_81#_c_2049_n 0.00183434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_415_81#_c_2050_n 0.00290125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_Q_c_2193_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_127 VNB N_Q_c_2194_n 0.00178889f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_128 VNB N_Q_c_2195_n 0.00200996f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_129 VNB Q 0.0195094f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_130 VNB N_VGND_c_2260_n 0.0110567f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_131 VNB N_VGND_c_2261_n 0.0138371f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_132 VNB N_VGND_c_2262_n 0.00496478f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_133 VNB N_VGND_c_2263_n 0.00428891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2264_n 0.00497485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2265_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2266_n 0.0413125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2267_n 0.0676218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2268_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2269_n 0.0194685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2270_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2271_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2272_n 0.0605088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2273_n 0.0602754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2274_n 0.0428668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2275_n 0.0151727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2276_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2277_n 0.0168909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2278_n 0.00808418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2279_n 0.00481148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2280_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2281_n 0.0272142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2282_n 0.808255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_noxref_24_c_2403_n 0.0143966f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_154 VNB N_noxref_24_c_2404_n 0.00655627f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.935
cc_155 VNB N_noxref_24_c_2405_n 0.0026149f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_156 VPB N_A_27_74#_c_306_n 0.0534868f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_157 VPB N_A_27_74#_c_302_n 0.016494f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_158 VPB N_A_27_74#_c_308_n 0.0338402f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_159 VPB N_A_27_74#_c_309_n 0.0351167f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_160 VPB N_A_27_74#_c_310_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_161 VPB N_A_27_74#_c_311_n 0.00370424f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_162 VPB N_SCE_c_390_n 0.0264922f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_163 VPB N_SCE_c_391_n 0.0318721f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_164 VPB N_SCE_c_392_n 0.0231924f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_165 VPB N_SCE_c_393_n 0.0275749f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_166 VPB N_SCE_c_384_n 0.00782879f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_167 VPB N_SCE_c_385_n 0.0410982f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_168 VPB N_SCE_c_387_n 0.00295534f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_169 VPB N_SCE_c_389_n 0.00270951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_D_c_470_n 0.030204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_D_c_475_n 0.0220375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_SCD_c_520_n 0.0170214f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_173 VPB N_SCD_c_517_n 0.0506499f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_174 VPB SCD 0.00172059f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_175 VPB N_RESET_B_M1023_g 0.0125834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_RESET_B_c_569_n 0.021814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_RESET_B_c_570_n 0.0167099f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_178 VPB N_RESET_B_c_566_n 0.0106437f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_179 VPB N_RESET_B_M1041_g 0.00996849f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_180 VPB N_RESET_B_c_573_n 0.0149978f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_181 VPB N_RESET_B_c_574_n 0.0251375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_RESET_B_c_575_n 0.0204581f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_183 VPB N_RESET_B_c_576_n 0.00161953f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_184 VPB N_RESET_B_c_577_n 0.0213442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_RESET_B_c_578_n 0.00238517f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_186 VPB N_RESET_B_c_579_n 0.00204342f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB RESET_B 0.00336207f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_188 VPB N_RESET_B_c_581_n 0.0662647f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_189 VPB N_RESET_B_c_582_n 0.00233009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_RESET_B_c_583_n 0.0621565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_RESET_B_c_584_n 0.00478311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_RESET_B_c_585_n 0.0461401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_CLK_c_768_n 0.0297761f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_194 VPB N_A_1034_74#_c_844_n 0.0145296f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.01
cc_195 VPB N_A_1034_74#_c_845_n 0.0198309f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_196 VPB N_A_1034_74#_c_823_n 0.0141763f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_197 VPB N_A_1034_74#_c_847_n 0.057308f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_198 VPB N_A_1034_74#_c_832_n 0.00168243f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_199 VPB N_A_1034_74#_c_837_n 0.00112381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1034_74#_c_850_n 0.00501177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1034_74#_c_839_n 0.00732078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1034_74#_c_843_n 0.0202793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_1367_112#_c_1048_n 0.0136749f $X=-0.19 $Y=1.66 $X2=2.495
+ $Y2=2.245
cc_204 VPB N_A_1367_112#_c_1049_n 0.0212139f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_205 VPB N_A_1367_112#_c_1044_n 0.00199812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1367_112#_c_1045_n 0.0360196f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_207 VPB N_A_1367_112#_c_1047_n 7.08723e-19 $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_208 VPB N_A_1367_112#_c_1053_n 0.00336227f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_209 VPB N_A_1233_138#_c_1153_n 0.0157054f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_210 VPB N_A_1233_138#_c_1161_n 0.0155175f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_211 VPB N_A_1233_138#_c_1162_n 0.0030701f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_212 VPB N_A_1233_138#_c_1154_n 0.00749326f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_213 VPB N_A_1233_138#_c_1155_n 0.0121924f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_214 VPB N_A_1233_138#_c_1158_n 0.00783535f $X=-0.19 $Y=1.66 $X2=2.54
+ $Y2=1.995
cc_215 VPB N_A_1233_138#_c_1166_n 0.00186797f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_855_368#_c_1288_n 0.0223719f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_217 VPB N_A_855_368#_c_1290_n 0.076923f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_218 VPB N_A_855_368#_c_1303_n 0.0586461f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_219 VPB N_A_855_368#_c_1304_n 0.0123764f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_220 VPB N_A_855_368#_c_1305_n 0.00718351f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_855_368#_c_1306_n 0.0163876f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_222 VPB N_A_855_368#_c_1307_n 0.0162442f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_223 VPB N_A_855_368#_c_1308_n 0.186352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_855_368#_c_1309_n 0.00735052f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_225 VPB N_A_855_368#_c_1310_n 0.0131075f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_226 VPB N_A_855_368#_M1003_g 0.0082806f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_227 VPB N_A_855_368#_c_1293_n 0.0195614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_855_368#_c_1294_n 0.00360844f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_229 VPB N_A_855_368#_c_1314_n 0.0089864f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_230 VPB N_A_855_368#_c_1315_n 0.00254706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_855_368#_c_1299_n 0.00276966f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_855_368#_c_1317_n 0.0018583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_2003_48#_c_1485_n 0.0412197f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_234 VPB N_A_2003_48#_c_1494_n 0.0232955f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_235 VPB N_A_2003_48#_c_1495_n 0.00836779f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_236 VPB N_A_2003_48#_c_1491_n 0.0185734f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_237 VPB N_A_1745_74#_c_1574_n 3.48694e-19 $X=-0.19 $Y=1.66 $X2=2.495
+ $Y2=2.245
cc_238 VPB N_A_1745_74#_c_1589_n 0.0451105f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_239 VPB N_A_1745_74#_c_1590_n 0.0242804f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_240 VPB N_A_1745_74#_c_1591_n 0.0157526f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_241 VPB N_A_1745_74#_c_1578_n 0.0115338f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_242 VPB N_A_1745_74#_c_1593_n 0.0157765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1745_74#_c_1580_n 0.00496747f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_244 VPB N_A_1745_74#_c_1595_n 0.00176961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1745_74#_c_1583_n 0.00118746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1745_74#_c_1597_n 0.0080022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1745_74#_c_1598_n 0.00237571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1745_74#_c_1599_n 0.00700686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_2339_74#_c_1748_n 0.0160879f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.935
cc_250 VPB N_A_2339_74#_c_1749_n 0.0148316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_2339_74#_c_1750_n 0.0143946f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_252 VPB N_A_2339_74#_c_1751_n 0.0165543f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_253 VPB N_A_2339_74#_c_1744_n 0.00394633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_2339_74#_c_1747_n 0.0271172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1855_n 0.0066125f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_256 VPB N_VPWR_c_1856_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1857_n 0.013846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1858_n 0.0230775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1859_n 0.0142717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1860_n 0.0137486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1861_n 0.0277893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1862_n 0.0214037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1863_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1864_n 0.00508939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1865_n 0.0115177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1866_n 0.0443867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1867_n 0.0375576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1868_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1869_n 0.0520927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1870_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1871_n 0.0191816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1872_n 0.0457766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1873_n 0.0618141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1874_n 0.0245819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1875_n 0.0218508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1876_n 0.0173667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1877_n 0.0312859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1878_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1879_n 0.00463502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1880_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1881_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1882_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1883_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1854_n 0.136739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_415_81#_c_2046_n 0.00482108f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_286 VPB N_A_415_81#_c_2052_n 0.00940845f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_287 VPB N_A_415_81#_c_2053_n 0.0125416f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_288 VPB N_A_415_81#_c_2054_n 0.00122623f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_289 VPB N_A_415_81#_c_2055_n 0.00722066f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_290 VPB N_A_415_81#_c_2050_n 0.00581282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_A_415_81#_c_2057_n 0.00257025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_A_415_81#_c_2058_n 0.00910856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_Q_c_2197_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_294 VPB N_Q_c_2198_n 0.0023624f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_295 VPB N_Q_c_2199_n 0.00183442f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_296 VPB N_Q_c_2200_n 0.00221952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB Q 0.0136248f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_298 N_A_27_74#_c_309_n N_SCE_c_390_n 0.0121883f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_310_n N_SCE_c_390_n 0.00496169f $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_301_n N_SCE_M1037_g 0.00686809f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_302_n N_SCE_M1037_g 0.00830473f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_303_n N_SCE_M1037_g 0.0281157f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_305_n N_SCE_M1037_g 0.0181297f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_308_n N_SCE_c_391_n 0.0173713f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_309_n N_SCE_c_391_n 0.00721429f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_310_n N_SCE_c_391_n 4.59028e-19 $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_309_n N_SCE_c_392_n 0.0100663f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_309_n N_SCE_c_393_n 0.00784761f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_306_n N_SCE_c_382_n 0.0165639f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_311_n N_SCE_c_382_n 3.28396e-19 $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_302_n N_SCE_c_384_n 0.0158921f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_303_n N_SCE_c_384_n 0.00162366f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_299_n N_SCE_c_385_n 0.0106974f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_303_n N_SCE_c_385_n 0.00180358f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_309_n N_SCE_c_385_n 0.0170396f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_305_n N_SCE_c_385_n 0.0175645f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_306_n N_SCE_c_386_n 2.04435e-19 $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_c_309_n N_SCE_c_386_n 0.0253562f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_311_n N_SCE_c_386_n 0.00219772f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_306_n N_SCE_c_387_n 0.00103776f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_321 N_A_27_74#_c_311_n N_SCE_c_387_n 0.0242605f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_299_n N_SCE_c_388_n 0.00818136f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_323 N_A_27_74#_c_302_n N_SCE_c_388_n 0.0170838f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_303_n N_SCE_c_388_n 0.0353374f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_325 N_A_27_74#_c_309_n N_SCE_c_388_n 0.0893268f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_326 N_A_27_74#_c_305_n N_SCE_c_388_n 0.00202099f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_306_n N_D_c_470_n 0.0183644f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_309_n N_D_c_470_n 0.00915555f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_311_n N_D_c_470_n 0.00125897f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_306_n N_D_c_475_n 0.0140909f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_309_n N_D_c_475_n 0.00753583f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_299_n N_D_c_471_n 0.00979811f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_333 N_A_27_74#_c_303_n N_D_c_471_n 2.46751e-19 $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_334 N_A_27_74#_c_305_n N_D_c_471_n 0.00223479f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_335 N_A_27_74#_c_300_n N_D_c_472_n 0.00580814f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_336 N_A_27_74#_c_303_n N_D_c_472_n 0.0143876f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_337 N_A_27_74#_c_305_n N_D_c_472_n 8.79717e-19 $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_338 N_A_27_74#_c_300_n N_D_c_473_n 0.0224455f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_339 N_A_27_74#_c_306_n N_SCD_c_520_n 0.0258628f $X=2.495 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_340 N_A_27_74#_c_306_n N_SCD_c_517_n 0.0203694f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_341 N_A_27_74#_c_311_n N_SCD_c_517_n 0.0015633f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_342 N_A_27_74#_c_306_n SCD 0.00117743f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_343 N_A_27_74#_c_311_n SCD 0.0182021f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_344 N_A_27_74#_c_306_n N_VPWR_c_1855_n 0.00141778f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_308_n N_VPWR_c_1871_n 0.0145938f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_306_n N_VPWR_c_1872_n 0.00445602f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_308_n N_VPWR_c_1877_n 0.0247088f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_309_n N_VPWR_c_1877_n 0.0746993f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_306_n N_VPWR_c_1854_n 0.00448781f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_308_n N_VPWR_c_1854_n 0.0120466f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_306_n N_A_415_81#_c_2059_n 0.010208f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_311_n N_A_415_81#_c_2059_n 0.0180834f $X=2.54 $Y=1.995 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_306_n N_A_415_81#_c_2057_n 0.00974144f $X=2.495 $Y=2.245
+ $X2=0 $Y2=0
cc_354 N_A_27_74#_c_309_n N_A_415_81#_c_2057_n 0.0189432f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_311_n N_A_415_81#_c_2057_n 0.00295889f $X=2.54 $Y=1.995
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_c_300_n N_VGND_c_2260_n 0.00287309f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_301_n N_VGND_c_2260_n 0.0156021f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_303_n N_VGND_c_2260_n 0.0254818f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_305_n N_VGND_c_2260_n 0.00149092f $X=0.975 $Y=1.01 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_300_n N_VGND_c_2267_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_301_n N_VGND_c_2271_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_301_n N_VGND_c_2282_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_300_n N_noxref_24_c_2403_n 0.011495f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_300_n N_noxref_24_c_2404_n 0.00899724f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_365 N_A_27_74#_c_303_n N_noxref_24_c_2404_n 0.00178881f $X=0.975 $Y=1.1 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_305_n N_noxref_24_c_2404_n 0.00859402f $X=0.975 $Y=1.01
+ $X2=0 $Y2=0
cc_367 N_SCE_c_385_n N_D_c_470_n 0.0203026f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_368 N_SCE_c_386_n N_D_c_470_n 0.0146397f $X=2.405 $Y=1.575 $X2=0 $Y2=0
cc_369 N_SCE_c_387_n N_D_c_470_n 3.21106e-19 $X=2.57 $Y=1.425 $X2=0 $Y2=0
cc_370 N_SCE_c_389_n N_D_c_470_n 0.00479409f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_371 N_SCE_c_392_n N_D_c_475_n 0.0203026f $X=1.625 $Y=2.155 $X2=0 $Y2=0
cc_372 N_SCE_c_393_n N_D_c_475_n 0.0373591f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_373 N_SCE_c_382_n N_D_c_471_n 0.0223603f $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_374 N_SCE_M1039_g N_D_c_471_n 0.00179056f $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_375 N_SCE_c_387_n N_D_c_471_n 0.00148517f $X=2.57 $Y=1.425 $X2=0 $Y2=0
cc_376 N_SCE_c_389_n N_D_c_471_n 0.00411836f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_377 N_SCE_c_382_n N_D_c_472_n 9.75781e-19 $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_378 N_SCE_M1039_g N_D_c_472_n 4.78719e-19 $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_379 N_SCE_c_385_n N_D_c_472_n 0.00106377f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_380 N_SCE_c_388_n N_D_c_472_n 0.0344941f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_381 N_SCE_M1039_g N_D_c_473_n 0.00976046f $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_382 N_SCE_c_382_n N_SCD_M1040_g 0.00891165f $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_383 N_SCE_M1039_g N_SCD_M1040_g 0.0494943f $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_384 N_SCE_c_387_n N_SCD_M1040_g 0.00105653f $X=2.57 $Y=1.425 $X2=0 $Y2=0
cc_385 N_SCE_c_382_n SCD 5.22436e-19 $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_386 N_SCE_c_387_n SCD 0.0142044f $X=2.57 $Y=1.425 $X2=0 $Y2=0
cc_387 N_SCE_c_382_n N_SCD_c_519_n 0.00914109f $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_388 N_SCE_c_387_n N_SCD_c_519_n 0.00206001f $X=2.57 $Y=1.425 $X2=0 $Y2=0
cc_389 N_SCE_c_391_n N_VPWR_c_1871_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_390 N_SCE_c_393_n N_VPWR_c_1872_n 0.00415318f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_391 N_SCE_c_391_n N_VPWR_c_1877_n 0.017697f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_392 N_SCE_c_393_n N_VPWR_c_1877_n 0.0163904f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_393 N_SCE_c_391_n N_VPWR_c_1854_n 0.00865213f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_394 N_SCE_c_393_n N_VPWR_c_1854_n 0.00817532f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_395 N_SCE_c_382_n N_A_415_81#_c_2044_n 0.00694815f $X=2.785 $Y=1.05 $X2=0
+ $Y2=0
cc_396 N_SCE_M1039_g N_A_415_81#_c_2044_n 0.0128765f $X=2.785 $Y=0.615 $X2=0
+ $Y2=0
cc_397 N_SCE_c_386_n N_A_415_81#_c_2044_n 0.00413271f $X=2.405 $Y=1.575 $X2=0
+ $Y2=0
cc_398 N_SCE_c_387_n N_A_415_81#_c_2044_n 0.019844f $X=2.57 $Y=1.425 $X2=0 $Y2=0
cc_399 N_SCE_c_382_n N_A_415_81#_c_2045_n 0.00571982f $X=2.785 $Y=1.05 $X2=0
+ $Y2=0
cc_400 N_SCE_M1039_g N_A_415_81#_c_2045_n 0.00628407f $X=2.785 $Y=0.615 $X2=0
+ $Y2=0
cc_401 N_SCE_c_393_n N_A_415_81#_c_2057_n 0.00182961f $X=1.625 $Y=2.245 $X2=0
+ $Y2=0
cc_402 N_SCE_M1037_g N_VGND_c_2260_n 0.0129468f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_403 N_SCE_M1039_g N_VGND_c_2267_n 9.15902e-19 $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_404 N_SCE_M1037_g N_VGND_c_2271_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_405 N_SCE_M1037_g N_VGND_c_2282_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_406 N_SCE_c_382_n N_noxref_24_c_2403_n 2.94195e-19 $X=2.785 $Y=1.05 $X2=0
+ $Y2=0
cc_407 N_SCE_M1039_g N_noxref_24_c_2403_n 0.0121157f $X=2.785 $Y=0.615 $X2=0
+ $Y2=0
cc_408 N_SCE_M1037_g N_noxref_24_c_2404_n 9.19966e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_409 N_SCE_M1039_g N_noxref_24_c_2405_n 0.00135222f $X=2.785 $Y=0.615 $X2=0
+ $Y2=0
cc_410 N_D_c_475_n N_VPWR_c_1872_n 0.00445602f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_411 N_D_c_475_n N_VPWR_c_1877_n 0.00236192f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_412 N_D_c_475_n N_VPWR_c_1854_n 0.00858241f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_413 N_D_c_471_n N_A_415_81#_c_2044_n 0.00121993f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_414 N_D_c_472_n N_A_415_81#_c_2044_n 0.0115884f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_415 N_D_c_473_n N_A_415_81#_c_2044_n 0.00599383f $X=1.952 $Y=0.935 $X2=0
+ $Y2=0
cc_416 N_D_c_475_n N_A_415_81#_c_2057_n 0.0112736f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_417 N_D_c_473_n N_VGND_c_2267_n 9.15902e-19 $X=1.952 $Y=0.935 $X2=0 $Y2=0
cc_418 N_D_c_471_n N_noxref_24_c_2403_n 0.00121903f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_419 N_D_c_472_n N_noxref_24_c_2403_n 0.014028f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_420 N_D_c_473_n N_noxref_24_c_2403_n 0.0125454f $X=1.952 $Y=0.935 $X2=0 $Y2=0
cc_421 N_D_c_473_n N_noxref_24_c_2404_n 0.00108287f $X=1.952 $Y=0.935 $X2=0
+ $Y2=0
cc_422 N_D_c_472_n noxref_25 0.00395662f $X=1.935 $Y=1.1 $X2=-0.19 $Y2=-0.245
cc_423 N_SCD_M1040_g N_RESET_B_M1023_g 0.0358944f $X=3.175 $Y=0.615 $X2=0 $Y2=0
cc_424 SCD N_RESET_B_M1023_g 4.27105e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_425 N_SCD_c_519_n N_RESET_B_M1023_g 0.0188651f $X=3.11 $Y=1.605 $X2=0 $Y2=0
cc_426 N_SCD_c_520_n N_RESET_B_c_569_n 0.0163026f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_427 N_SCD_c_517_n N_RESET_B_c_581_n 0.018487f $X=3.11 $Y=1.945 $X2=0 $Y2=0
cc_428 SCD N_RESET_B_c_581_n 4.34698e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_429 N_SCD_c_520_n N_VPWR_c_1855_n 0.0100582f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_430 N_SCD_c_520_n N_VPWR_c_1872_n 0.00413917f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_431 N_SCD_c_520_n N_VPWR_c_1854_n 0.00409681f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_432 N_SCD_M1040_g N_A_415_81#_c_2044_n 0.00137126f $X=3.175 $Y=0.615 $X2=0
+ $Y2=0
cc_433 N_SCD_c_520_n N_A_415_81#_c_2059_n 0.0130079f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_434 N_SCD_c_517_n N_A_415_81#_c_2059_n 8.17297e-19 $X=3.11 $Y=1.945 $X2=0
+ $Y2=0
cc_435 SCD N_A_415_81#_c_2059_n 0.0212424f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_436 N_SCD_M1040_g N_A_415_81#_c_2045_n 0.0124697f $X=3.175 $Y=0.615 $X2=0
+ $Y2=0
cc_437 SCD N_A_415_81#_c_2045_n 0.0146824f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_438 N_SCD_c_519_n N_A_415_81#_c_2045_n 0.00106346f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_439 N_SCD_c_520_n N_A_415_81#_c_2046_n 0.00151656f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_440 N_SCD_M1040_g N_A_415_81#_c_2046_n 0.0070009f $X=3.175 $Y=0.615 $X2=0
+ $Y2=0
cc_441 N_SCD_c_517_n N_A_415_81#_c_2046_n 0.00183512f $X=3.11 $Y=1.945 $X2=0
+ $Y2=0
cc_442 SCD N_A_415_81#_c_2046_n 0.0534507f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_443 N_SCD_c_519_n N_A_415_81#_c_2046_n 0.0038704f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_444 N_SCD_c_520_n N_A_415_81#_c_2052_n 4.52461e-19 $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_445 N_SCD_c_520_n N_A_415_81#_c_2054_n 5.56969e-19 $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_446 N_SCD_c_520_n N_A_415_81#_c_2057_n 0.00167919f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_447 N_SCD_M1040_g N_VGND_c_2267_n 9.09582e-19 $X=3.175 $Y=0.615 $X2=0 $Y2=0
cc_448 N_SCD_M1040_g N_noxref_24_c_2403_n 0.00856921f $X=3.175 $Y=0.615 $X2=0
+ $Y2=0
cc_449 N_SCD_M1040_g N_noxref_24_c_2405_n 0.00853984f $X=3.175 $Y=0.615 $X2=0
+ $Y2=0
cc_450 N_RESET_B_c_575_n N_CLK_c_768_n 0.00217884f $X=7.775 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_451 N_RESET_B_c_581_n N_CLK_c_768_n 0.00390967f $X=3.605 $Y=2.037 $X2=-0.19
+ $Y2=-0.245
cc_452 N_RESET_B_c_582_n N_CLK_c_768_n 4.10166e-19 $X=3.95 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_453 N_RESET_B_M1023_g N_CLK_c_770_n 0.013532f $X=3.605 $Y=0.615 $X2=0 $Y2=0
cc_454 N_RESET_B_c_575_n N_CLK_c_770_n 0.00236558f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_455 N_RESET_B_c_576_n N_CLK_c_770_n 0.00141283f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_456 N_RESET_B_c_581_n N_CLK_c_770_n 0.00776499f $X=3.605 $Y=2.037 $X2=0 $Y2=0
cc_457 N_RESET_B_c_582_n N_CLK_c_770_n 0.00164317f $X=3.95 $Y=1.995 $X2=0 $Y2=0
cc_458 N_RESET_B_c_575_n N_CLK_c_781_n 0.0055638f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_459 N_RESET_B_M1023_g N_CLK_c_771_n 0.00261733f $X=3.605 $Y=0.615 $X2=0 $Y2=0
cc_460 N_RESET_B_c_576_n N_CLK_c_771_n 0.003583f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_461 N_RESET_B_c_581_n N_CLK_c_771_n 5.51696e-19 $X=3.605 $Y=2.037 $X2=0 $Y2=0
cc_462 N_RESET_B_c_582_n N_CLK_c_771_n 0.0104506f $X=3.95 $Y=1.995 $X2=0 $Y2=0
cc_463 N_RESET_B_c_575_n N_A_1034_74#_c_844_n 0.003934f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_464 N_RESET_B_c_575_n N_A_1034_74#_c_823_n 0.00392629f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_465 N_RESET_B_c_577_n N_A_1034_74#_c_847_n 0.00245933f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_466 N_RESET_B_c_575_n N_A_1034_74#_c_832_n 0.0168899f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_467 N_RESET_B_c_563_n N_A_1034_74#_c_833_n 0.0104f $X=7.3 $Y=1.185 $X2=0
+ $Y2=0
cc_468 N_RESET_B_c_563_n N_A_1034_74#_c_858_n 4.46705e-19 $X=7.3 $Y=1.185 $X2=0
+ $Y2=0
cc_469 N_RESET_B_c_577_n N_A_1034_74#_c_837_n 0.0104861f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_470 N_RESET_B_c_577_n N_A_1034_74#_c_860_n 0.00467739f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_471 N_RESET_B_c_577_n N_A_1034_74#_c_850_n 0.0172592f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_472 N_RESET_B_c_575_n N_A_1034_74#_c_839_n 0.0309583f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_473 N_RESET_B_c_563_n N_A_1034_74#_c_840_n 0.00237513f $X=7.3 $Y=1.185 $X2=0
+ $Y2=0
cc_474 N_RESET_B_c_575_n N_A_1034_74#_c_843_n 0.00388711f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_475 N_RESET_B_c_563_n N_A_1367_112#_M1001_g 0.0394201f $X=7.3 $Y=1.185 $X2=0
+ $Y2=0
cc_476 N_RESET_B_c_566_n N_A_1367_112#_M1001_g 0.00326496f $X=7.67 $Y=1.82 $X2=0
+ $Y2=0
cc_477 N_RESET_B_c_575_n N_A_1367_112#_c_1048_n 0.0105234f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_478 N_RESET_B_c_583_n N_A_1367_112#_c_1048_n 0.00683215f $X=7.67 $Y=2.03
+ $X2=0 $Y2=0
cc_479 N_RESET_B_c_570_n N_A_1367_112#_c_1049_n 0.0123322f $X=7.665 $Y=2.24
+ $X2=0 $Y2=0
cc_480 N_RESET_B_c_563_n N_A_1367_112#_c_1044_n 0.00515512f $X=7.3 $Y=1.185
+ $X2=0 $Y2=0
cc_481 N_RESET_B_c_565_n N_A_1367_112#_c_1044_n 0.00753567f $X=7.375 $Y=1.26
+ $X2=0 $Y2=0
cc_482 N_RESET_B_c_566_n N_A_1367_112#_c_1044_n 0.00113842f $X=7.67 $Y=1.82
+ $X2=0 $Y2=0
cc_483 N_RESET_B_c_575_n N_A_1367_112#_c_1044_n 0.009228f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_484 N_RESET_B_c_565_n N_A_1367_112#_c_1045_n 0.00620241f $X=7.375 $Y=1.26
+ $X2=0 $Y2=0
cc_485 N_RESET_B_c_566_n N_A_1367_112#_c_1045_n 0.0110407f $X=7.67 $Y=1.82 $X2=0
+ $Y2=0
cc_486 N_RESET_B_c_575_n N_A_1367_112#_c_1045_n 0.00237054f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_487 N_RESET_B_c_583_n N_A_1367_112#_c_1045_n 0.00760267f $X=7.67 $Y=2.03
+ $X2=0 $Y2=0
cc_488 N_RESET_B_c_563_n N_A_1367_112#_c_1067_n 0.00422682f $X=7.3 $Y=1.185
+ $X2=0 $Y2=0
cc_489 N_RESET_B_c_577_n N_A_1367_112#_c_1047_n 0.00727956f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_490 N_RESET_B_c_577_n N_A_1367_112#_c_1053_n 0.030687f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_491 N_RESET_B_c_563_n N_A_1367_112#_c_1070_n 0.0067801f $X=7.3 $Y=1.185 $X2=0
+ $Y2=0
cc_492 N_RESET_B_c_564_n N_A_1367_112#_c_1070_n 0.00975109f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_493 N_RESET_B_c_564_n N_A_1233_138#_M1025_g 0.00269339f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_494 N_RESET_B_c_577_n N_A_1233_138#_c_1153_n 3.01246e-19 $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_495 N_RESET_B_c_577_n N_A_1233_138#_c_1161_n 0.00699288f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_496 N_RESET_B_c_575_n N_A_1233_138#_c_1162_n 0.00819966f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_497 N_RESET_B_c_563_n N_A_1233_138#_c_1171_n 2.03434e-19 $X=7.3 $Y=1.185
+ $X2=0 $Y2=0
cc_498 N_RESET_B_c_563_n N_A_1233_138#_c_1154_n 2.11405e-19 $X=7.3 $Y=1.185
+ $X2=0 $Y2=0
cc_499 N_RESET_B_c_575_n N_A_1233_138#_c_1154_n 0.0241128f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_500 N_RESET_B_c_575_n N_A_1233_138#_c_1174_n 0.020887f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_501 N_RESET_B_c_570_n N_A_1233_138#_c_1155_n 0.0179696f $X=7.665 $Y=2.24
+ $X2=0 $Y2=0
cc_502 N_RESET_B_c_566_n N_A_1233_138#_c_1155_n 0.0117416f $X=7.67 $Y=1.82 $X2=0
+ $Y2=0
cc_503 N_RESET_B_c_575_n N_A_1233_138#_c_1155_n 0.0257004f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_504 N_RESET_B_c_578_n N_A_1233_138#_c_1155_n 0.0106292f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_505 N_RESET_B_c_579_n N_A_1233_138#_c_1155_n 0.0363198f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_506 N_RESET_B_c_583_n N_A_1233_138#_c_1155_n 0.020253f $X=7.67 $Y=2.03 $X2=0
+ $Y2=0
cc_507 N_RESET_B_c_564_n N_A_1233_138#_c_1156_n 0.00569114f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_508 N_RESET_B_c_566_n N_A_1233_138#_c_1156_n 0.00438308f $X=7.67 $Y=1.82
+ $X2=0 $Y2=0
cc_509 N_RESET_B_c_564_n N_A_1233_138#_c_1157_n 0.00188178f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_510 N_RESET_B_c_566_n N_A_1233_138#_c_1157_n 0.00586797f $X=7.67 $Y=1.82
+ $X2=0 $Y2=0
cc_511 N_RESET_B_c_575_n N_A_1233_138#_c_1157_n 0.00357593f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_512 N_RESET_B_c_577_n N_A_1233_138#_c_1157_n 0.00641796f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_513 N_RESET_B_c_578_n N_A_1233_138#_c_1157_n 0.00373314f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_514 N_RESET_B_c_579_n N_A_1233_138#_c_1157_n 0.0158779f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_515 N_RESET_B_c_583_n N_A_1233_138#_c_1157_n 0.00716371f $X=7.67 $Y=2.03
+ $X2=0 $Y2=0
cc_516 N_RESET_B_c_564_n N_A_1233_138#_c_1158_n 0.0194698f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_517 N_RESET_B_c_577_n N_A_1233_138#_c_1158_n 0.00591166f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_518 N_RESET_B_c_579_n N_A_1233_138#_c_1158_n 6.12607e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_519 N_RESET_B_c_583_n N_A_1233_138#_c_1158_n 0.00918526f $X=7.67 $Y=2.03
+ $X2=0 $Y2=0
cc_520 N_RESET_B_c_575_n N_A_855_368#_M1019_s 0.0011702f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_521 N_RESET_B_c_575_n N_A_855_368#_c_1288_n 0.00496452f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_522 N_RESET_B_c_575_n N_A_855_368#_c_1290_n 0.00533173f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_523 N_RESET_B_c_575_n N_A_855_368#_c_1307_n 0.00397216f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_524 N_RESET_B_c_570_n N_A_855_368#_c_1308_n 0.0100134f $X=7.665 $Y=2.24 $X2=0
+ $Y2=0
cc_525 N_RESET_B_c_577_n N_A_855_368#_M1003_g 0.0124871f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_526 N_RESET_B_c_577_n N_A_855_368#_c_1293_n 0.00423021f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_527 N_RESET_B_M1023_g N_A_855_368#_c_1297_n 0.00403112f $X=3.605 $Y=0.615
+ $X2=0 $Y2=0
cc_528 N_RESET_B_M1023_g N_A_855_368#_c_1326_n 0.00402378f $X=3.605 $Y=0.615
+ $X2=0 $Y2=0
cc_529 N_RESET_B_c_575_n N_A_855_368#_c_1315_n 0.0157342f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_530 N_RESET_B_M1023_g N_A_855_368#_c_1317_n 2.07062e-19 $X=3.605 $Y=0.615
+ $X2=0 $Y2=0
cc_531 N_RESET_B_c_575_n N_A_855_368#_c_1317_n 0.014404f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_532 N_RESET_B_c_576_n N_A_855_368#_c_1317_n 0.00277564f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_581_n N_A_855_368#_c_1317_n 0.0023658f $X=3.605 $Y=2.037
+ $X2=0 $Y2=0
cc_534 N_RESET_B_c_582_n N_A_855_368#_c_1317_n 0.0240037f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_575_n N_A_855_368#_c_1300_n 0.00697206f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_536 N_RESET_B_M1041_g N_A_2003_48#_M1028_g 0.0216011f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_537 N_RESET_B_c_573_n N_A_2003_48#_c_1485_n 0.00394367f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_577_n N_A_2003_48#_c_1485_n 0.00331802f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_584_n N_A_2003_48#_c_1485_n 0.00106389f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_540 N_RESET_B_c_585_n N_A_2003_48#_c_1485_n 0.029932f $X=10.94 $Y=1.985 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_574_n N_A_2003_48#_c_1494_n 0.0126655f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_542 N_RESET_B_M1041_g N_A_2003_48#_c_1486_n 0.0128807f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_577_n N_A_2003_48#_c_1486_n 0.00879069f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_544 RESET_B N_A_2003_48#_c_1486_n 0.00259932f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_545 N_RESET_B_c_584_n N_A_2003_48#_c_1486_n 0.0152297f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_585_n N_A_2003_48#_c_1486_n 0.00391331f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_547 N_RESET_B_M1041_g N_A_2003_48#_c_1487_n 9.6789e-19 $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_548 N_RESET_B_M1041_g N_A_2003_48#_c_1489_n 0.00118187f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_549 N_RESET_B_c_577_n N_A_2003_48#_c_1489_n 0.00250381f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_550 N_RESET_B_M1041_g N_A_2003_48#_c_1490_n 0.029932f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_551 N_RESET_B_c_574_n N_A_2003_48#_c_1495_n 0.00739105f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_552 N_RESET_B_M1041_g N_A_2003_48#_c_1491_n 0.00453304f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_553 N_RESET_B_c_574_n N_A_2003_48#_c_1491_n 0.00121218f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_554 RESET_B N_A_2003_48#_c_1491_n 0.00621393f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_555 N_RESET_B_c_584_n N_A_2003_48#_c_1491_n 0.0154382f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_556 N_RESET_B_c_585_n N_A_2003_48#_c_1491_n 0.0101596f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_557 N_RESET_B_c_577_n N_A_1745_74#_M1003_d 0.00323029f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_558 N_RESET_B_M1041_g N_A_1745_74#_c_1573_n 0.0694909f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_585_n N_A_1745_74#_c_1589_n 0.00857472f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_560 N_RESET_B_c_573_n N_A_1745_74#_c_1590_n 0.00857472f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_574_n N_A_1745_74#_c_1590_n 0.010499f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_562 N_RESET_B_M1041_g N_A_1745_74#_c_1579_n 0.00550286f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_563 N_RESET_B_c_577_n N_A_1745_74#_c_1595_n 0.00708586f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_564 N_RESET_B_M1041_g N_A_1745_74#_c_1584_n 0.0150978f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_565 N_RESET_B_M1041_g N_A_1745_74#_c_1597_n 8.1654e-19 $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_577_n N_A_1745_74#_c_1597_n 0.0117357f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_567 N_RESET_B_c_584_n N_A_1745_74#_c_1597_n 0.00391217f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_568 N_RESET_B_c_577_n N_A_1745_74#_c_1598_n 0.00499654f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_569 N_RESET_B_c_573_n N_A_1745_74#_c_1599_n 0.00158772f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_570 N_RESET_B_c_574_n N_A_1745_74#_c_1599_n 2.73747e-19 $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_571 N_RESET_B_c_577_n N_A_1745_74#_c_1599_n 0.0200435f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_572 RESET_B N_A_1745_74#_c_1599_n 4.97327e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_573 N_RESET_B_c_584_n N_A_1745_74#_c_1599_n 0.00972451f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_585_n N_A_1745_74#_c_1599_n 8.72425e-19 $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_575 N_RESET_B_M1041_g N_A_1745_74#_c_1586_n 0.00118187f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_576 N_RESET_B_c_585_n N_A_1745_74#_c_1587_n 0.00231637f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_577 N_RESET_B_c_575_n N_VPWR_M1019_d 0.00316858f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_577_n N_VPWR_M1000_s 0.00641842f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_579 N_RESET_B_c_569_n N_VPWR_c_1855_n 0.00548967f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_580 N_RESET_B_c_570_n N_VPWR_c_1857_n 0.00421039f $X=7.665 $Y=2.24 $X2=0
+ $Y2=0
cc_581 N_RESET_B_c_575_n N_VPWR_c_1857_n 7.46496e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_570_n N_VPWR_c_1859_n 0.00486917f $X=7.665 $Y=2.24 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_566_n N_VPWR_c_1859_n 0.00160044f $X=7.67 $Y=1.82 $X2=0 $Y2=0
cc_584 N_RESET_B_c_577_n N_VPWR_c_1859_n 0.0183166f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_585 N_RESET_B_c_578_n N_VPWR_c_1859_n 5.40997e-19 $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_579_n N_VPWR_c_1859_n 0.0179605f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_587 N_RESET_B_c_583_n N_VPWR_c_1859_n 0.00312179f $X=7.67 $Y=2.03 $X2=0 $Y2=0
cc_588 N_RESET_B_c_574_n N_VPWR_c_1860_n 0.00816134f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_589 N_RESET_B_c_577_n N_VPWR_c_1860_n 0.00540169f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_590 RESET_B N_VPWR_c_1860_n 0.00113612f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_591 N_RESET_B_c_584_n N_VPWR_c_1860_n 0.00684931f $X=10.75 $Y=1.985 $X2=0
+ $Y2=0
cc_592 N_RESET_B_c_585_n N_VPWR_c_1860_n 0.00269311f $X=10.94 $Y=1.985 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_569_n N_VPWR_c_1867_n 0.00388952f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_594 N_RESET_B_c_574_n N_VPWR_c_1874_n 0.00445602f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_595 N_RESET_B_c_569_n N_VPWR_c_1854_n 0.00420469f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_570_n N_VPWR_c_1854_n 9.39239e-19 $X=7.665 $Y=2.24 $X2=0
+ $Y2=0
cc_597 N_RESET_B_c_574_n N_VPWR_c_1854_n 0.0089746f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_598 N_RESET_B_M1023_g N_A_415_81#_c_2045_n 0.0142027f $X=3.605 $Y=0.615 $X2=0
+ $Y2=0
cc_599 N_RESET_B_M1023_g N_A_415_81#_c_2046_n 0.0263717f $X=3.605 $Y=0.615 $X2=0
+ $Y2=0
cc_600 N_RESET_B_c_569_n N_A_415_81#_c_2046_n 0.00445911f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_601 N_RESET_B_c_576_n N_A_415_81#_c_2046_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_602 N_RESET_B_c_581_n N_A_415_81#_c_2046_n 0.0143328f $X=3.605 $Y=2.037 $X2=0
+ $Y2=0
cc_603 N_RESET_B_c_582_n N_A_415_81#_c_2046_n 0.0228135f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_604 N_RESET_B_c_569_n N_A_415_81#_c_2052_n 0.00791994f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_605 N_RESET_B_c_575_n N_A_415_81#_c_2053_n 0.0293302f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_606 N_RESET_B_c_576_n N_A_415_81#_c_2053_n 0.00388056f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_RESET_B_c_581_n N_A_415_81#_c_2053_n 0.00258186f $X=3.605 $Y=2.037
+ $X2=0 $Y2=0
cc_608 N_RESET_B_c_582_n N_A_415_81#_c_2053_n 0.00903824f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_569_n N_A_415_81#_c_2054_n 0.0119912f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_610 N_RESET_B_c_576_n N_A_415_81#_c_2054_n 4.98701e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_611 N_RESET_B_c_581_n N_A_415_81#_c_2054_n 0.00783424f $X=3.605 $Y=2.037
+ $X2=0 $Y2=0
cc_612 N_RESET_B_c_582_n N_A_415_81#_c_2054_n 0.0168153f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_613 N_RESET_B_c_575_n N_A_415_81#_c_2048_n 0.00381691f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_614 N_RESET_B_c_575_n N_A_415_81#_c_2055_n 0.016125f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_615 N_RESET_B_c_575_n N_A_415_81#_c_2050_n 0.011933f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_575_n N_A_415_81#_c_2058_n 0.0203963f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_617 N_RESET_B_M1023_g N_VGND_c_2261_n 0.00962592f $X=3.605 $Y=0.615 $X2=0
+ $Y2=0
cc_618 N_RESET_B_M1041_g N_VGND_c_2263_n 0.0101056f $X=10.63 $Y=0.58 $X2=0 $Y2=0
cc_619 N_RESET_B_M1023_g N_VGND_c_2267_n 0.00478603f $X=3.605 $Y=0.615 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_563_n N_VGND_c_2272_n 0.00294166f $X=7.3 $Y=1.185 $X2=0 $Y2=0
cc_621 N_RESET_B_M1041_g N_VGND_c_2274_n 0.00383152f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_622 N_RESET_B_M1023_g N_VGND_c_2282_n 0.0044912f $X=3.605 $Y=0.615 $X2=0
+ $Y2=0
cc_623 N_RESET_B_c_563_n N_VGND_c_2282_n 0.00451834f $X=7.3 $Y=1.185 $X2=0 $Y2=0
cc_624 N_RESET_B_M1041_g N_VGND_c_2282_n 0.0075694f $X=10.63 $Y=0.58 $X2=0 $Y2=0
cc_625 N_RESET_B_M1023_g N_noxref_24_c_2405_n 0.00724724f $X=3.605 $Y=0.615
+ $X2=0 $Y2=0
cc_626 N_CLK_M1007_g N_A_1034_74#_c_828_n 5.92939e-19 $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_627 N_CLK_c_768_n N_A_1034_74#_c_839_n 8.59843e-19 $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_628 N_CLK_M1007_g N_A_855_368#_c_1287_n 0.0228821f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_629 N_CLK_c_768_n N_A_855_368#_c_1288_n 0.048385f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_630 N_CLK_M1007_g N_A_855_368#_c_1288_n 0.0244578f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_631 N_CLK_c_781_n N_A_855_368#_c_1288_n 2.49644e-19 $X=4.47 $Y=1.425 $X2=0
+ $Y2=0
cc_632 N_CLK_M1007_g N_A_855_368#_c_1297_n 8.21824e-19 $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_633 N_CLK_M1007_g N_A_855_368#_c_1339_n 0.0148078f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_634 N_CLK_c_781_n N_A_855_368#_c_1339_n 0.00520588f $X=4.47 $Y=1.425 $X2=0
+ $Y2=0
cc_635 N_CLK_c_770_n N_A_855_368#_c_1326_n 0.00395112f $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_636 N_CLK_c_781_n N_A_855_368#_c_1326_n 0.0139041f $X=4.47 $Y=1.425 $X2=0
+ $Y2=0
cc_637 N_CLK_c_768_n N_A_855_368#_c_1315_n 0.0118317f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_638 N_CLK_c_781_n N_A_855_368#_c_1315_n 0.00251956f $X=4.47 $Y=1.425 $X2=0
+ $Y2=0
cc_639 N_CLK_M1007_g N_A_855_368#_c_1298_n 0.00285776f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_640 N_CLK_c_771_n N_A_855_368#_c_1298_n 0.00201078f $X=4.195 $Y=1.385 $X2=0
+ $Y2=0
cc_641 N_CLK_c_768_n N_A_855_368#_c_1299_n 0.00550019f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_642 N_CLK_c_781_n N_A_855_368#_c_1299_n 0.00111736f $X=4.47 $Y=1.425 $X2=0
+ $Y2=0
cc_643 N_CLK_c_768_n N_A_855_368#_c_1317_n 0.00541631f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_644 N_CLK_c_770_n N_A_855_368#_c_1317_n 0.004824f $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_645 N_CLK_c_781_n N_A_855_368#_c_1317_n 0.0144756f $X=4.47 $Y=1.425 $X2=0
+ $Y2=0
cc_646 N_CLK_M1007_g N_A_855_368#_c_1300_n 0.00271251f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_647 N_CLK_c_781_n N_A_855_368#_c_1300_n 0.0271023f $X=4.47 $Y=1.425 $X2=0
+ $Y2=0
cc_648 N_CLK_c_771_n N_A_855_368#_c_1300_n 4.76529e-19 $X=4.195 $Y=1.385 $X2=0
+ $Y2=0
cc_649 N_CLK_c_768_n N_VPWR_c_1856_n 0.0172823f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_650 N_CLK_c_768_n N_VPWR_c_1867_n 0.00413917f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_651 N_CLK_c_768_n N_VPWR_c_1854_n 0.00403443f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_652 N_CLK_c_770_n N_A_415_81#_c_2046_n 3.82626e-19 $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_653 N_CLK_c_771_n N_A_415_81#_c_2046_n 0.017388f $X=4.195 $Y=1.385 $X2=0
+ $Y2=0
cc_654 N_CLK_c_768_n N_A_415_81#_c_2052_n 0.0103912f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_655 N_CLK_c_768_n N_A_415_81#_c_2053_n 0.0146064f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_656 N_CLK_c_768_n N_A_415_81#_c_2054_n 0.00160388f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_657 N_CLK_M1007_g N_VGND_c_2261_n 0.00263389f $X=4.665 $Y=0.74 $X2=0 $Y2=0
cc_658 N_CLK_c_770_n N_VGND_c_2261_n 5.38625e-19 $X=4.555 $Y=1.425 $X2=0 $Y2=0
cc_659 N_CLK_c_771_n N_VGND_c_2261_n 0.00406664f $X=4.195 $Y=1.385 $X2=0 $Y2=0
cc_660 N_CLK_M1007_g N_VGND_c_2262_n 0.00883079f $X=4.665 $Y=0.74 $X2=0 $Y2=0
cc_661 N_CLK_M1007_g N_VGND_c_2269_n 0.00383152f $X=4.665 $Y=0.74 $X2=0 $Y2=0
cc_662 N_CLK_M1007_g N_VGND_c_2282_n 0.00762539f $X=4.665 $Y=0.74 $X2=0 $Y2=0
cc_663 N_A_1034_74#_c_834_n N_A_1367_112#_M1025_d 0.00224844f $X=8.825 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_664 N_A_1034_74#_M1016_g N_A_1367_112#_M1001_g 0.030435f $X=6.52 $Y=0.9 $X2=0
+ $Y2=0
cc_665 N_A_1034_74#_c_830_n N_A_1367_112#_M1001_g 0.00633573f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_666 N_A_1034_74#_c_840_n N_A_1367_112#_M1001_g 0.00342215f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_667 N_A_1034_74#_c_844_n N_A_1367_112#_c_1048_n 0.00142315f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_668 N_A_1034_74#_c_845_n N_A_1367_112#_c_1049_n 0.00142315f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_669 N_A_1034_74#_c_844_n N_A_1367_112#_c_1045_n 3.5795e-19 $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_670 N_A_1034_74#_c_823_n N_A_1367_112#_c_1045_n 0.030435f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_671 N_A_1034_74#_c_843_n N_A_1367_112#_c_1045_n 0.0023084f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_672 N_A_1034_74#_c_833_n N_A_1367_112#_c_1067_n 0.00761753f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_673 N_A_1034_74#_c_840_n N_A_1367_112#_c_1067_n 0.00974988f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_674 N_A_1034_74#_c_827_n N_A_1367_112#_c_1046_n 0.00476106f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_675 N_A_1034_74#_c_837_n N_A_1367_112#_c_1046_n 0.00539231f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_676 N_A_1034_74#_c_842_n N_A_1367_112#_c_1046_n 0.0108396f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_677 N_A_1034_74#_c_827_n N_A_1367_112#_c_1047_n 0.00855892f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_678 N_A_1034_74#_c_837_n N_A_1367_112#_c_1047_n 0.0129187f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_679 N_A_1034_74#_c_842_n N_A_1367_112#_c_1047_n 0.0180376f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_680 N_A_1034_74#_c_847_n N_A_1367_112#_c_1053_n 0.00106238f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_681 N_A_1034_74#_c_837_n N_A_1367_112#_c_1053_n 0.0240786f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_682 N_A_1034_74#_c_860_n N_A_1367_112#_c_1053_n 0.0118335f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_683 N_A_1034_74#_c_833_n N_A_1367_112#_c_1070_n 0.0484504f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_684 N_A_1034_74#_c_834_n N_A_1367_112#_c_1070_n 0.00422751f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_685 N_A_1034_74#_c_825_n N_A_1367_112#_c_1094_n 0.00932475f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_686 N_A_1034_74#_c_827_n N_A_1367_112#_c_1094_n 2.66567e-19 $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_687 N_A_1034_74#_c_834_n N_A_1367_112#_c_1094_n 0.02112f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_688 N_A_1034_74#_c_836_n N_A_1367_112#_c_1094_n 0.0232075f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_689 N_A_1034_74#_c_842_n N_A_1367_112#_c_1094_n 0.0158476f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_690 N_A_1034_74#_c_825_n N_A_1233_138#_M1025_g 0.0216734f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_691 N_A_1034_74#_c_833_n N_A_1233_138#_M1025_g 0.00459622f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_692 N_A_1034_74#_c_834_n N_A_1233_138#_M1025_g 0.00898149f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_693 N_A_1034_74#_c_835_n N_A_1233_138#_M1025_g 0.00298755f $X=8.1 $Y=0.34
+ $X2=0 $Y2=0
cc_694 N_A_1034_74#_c_827_n N_A_1233_138#_c_1153_n 0.0121912f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_695 N_A_1034_74#_c_837_n N_A_1233_138#_c_1153_n 3.24532e-19 $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_696 N_A_1034_74#_c_845_n N_A_1233_138#_c_1162_n 0.00181956f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_697 N_A_1034_74#_c_823_n N_A_1233_138#_c_1162_n 6.88374e-19 $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_698 N_A_1034_74#_M1016_g N_A_1233_138#_c_1171_n 0.00967614f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_699 N_A_1034_74#_c_830_n N_A_1233_138#_c_1171_n 0.0143872f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_700 N_A_1034_74#_c_844_n N_A_1233_138#_c_1154_n 3.69789e-19 $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_701 N_A_1034_74#_M1016_g N_A_1233_138#_c_1154_n 0.00659846f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_702 N_A_1034_74#_c_823_n N_A_1233_138#_c_1159_n 4.04338e-19 $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_703 N_A_1034_74#_M1016_g N_A_1233_138#_c_1159_n 0.0059346f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_704 N_A_1034_74#_c_830_n N_A_1233_138#_c_1159_n 0.0250791f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_705 N_A_1034_74#_c_840_n N_A_1233_138#_c_1159_n 0.00225536f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_706 N_A_1034_74#_c_828_n N_A_855_368#_c_1287_n 0.00431058f $X=5.31 $Y=0.515
+ $X2=0 $Y2=0
cc_707 N_A_1034_74#_c_829_n N_A_855_368#_c_1287_n 0.00186373f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_708 N_A_1034_74#_c_831_n N_A_855_368#_c_1287_n 0.00292953f $X=5.62 $Y=0.415
+ $X2=0 $Y2=0
cc_709 N_A_1034_74#_c_838_n N_A_855_368#_c_1287_n 0.00342133f $X=5.382 $Y=1.075
+ $X2=0 $Y2=0
cc_710 N_A_1034_74#_c_829_n N_A_855_368#_c_1288_n 7.82628e-19 $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_711 N_A_1034_74#_c_838_n N_A_855_368#_c_1288_n 0.0060592f $X=5.382 $Y=1.075
+ $X2=0 $Y2=0
cc_712 N_A_1034_74#_c_839_n N_A_855_368#_c_1288_n 0.0126368f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_713 N_A_1034_74#_c_829_n N_A_855_368#_c_1289_n 0.00601007f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_714 N_A_1034_74#_c_839_n N_A_855_368#_c_1289_n 0.00154346f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_715 N_A_1034_74#_c_844_n N_A_855_368#_c_1290_n 0.0108667f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_716 N_A_1034_74#_c_845_n N_A_855_368#_c_1290_n 0.0128837f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_717 N_A_1034_74#_c_829_n N_A_855_368#_c_1290_n 0.0104459f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_718 N_A_1034_74#_c_832_n N_A_855_368#_c_1290_n 0.0096323f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_719 N_A_1034_74#_c_839_n N_A_855_368#_c_1290_n 0.013478f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_720 N_A_1034_74#_c_843_n N_A_855_368#_c_1290_n 0.0213768f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_721 N_A_1034_74#_c_830_n N_A_855_368#_c_1291_n 3.42565e-19 $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_722 N_A_1034_74#_c_832_n N_A_855_368#_c_1291_n 0.00440403f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_723 N_A_1034_74#_c_843_n N_A_855_368#_c_1291_n 0.0143556f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_724 N_A_1034_74#_c_845_n N_A_855_368#_c_1303_n 0.0103487f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_725 N_A_1034_74#_M1016_g N_A_855_368#_c_1292_n 0.0189685f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_726 N_A_1034_74#_c_828_n N_A_855_368#_c_1292_n 0.00427211f $X=5.31 $Y=0.515
+ $X2=0 $Y2=0
cc_727 N_A_1034_74#_c_830_n N_A_855_368#_c_1292_n 0.00661564f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_728 N_A_1034_74#_c_845_n N_A_855_368#_c_1305_n 0.0024093f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_729 N_A_1034_74#_c_845_n N_A_855_368#_c_1307_n 0.0137651f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_730 N_A_1034_74#_c_823_n N_A_855_368#_c_1307_n 0.00110708f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_731 N_A_1034_74#_c_847_n N_A_855_368#_c_1309_n 0.00689629f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_732 N_A_1034_74#_c_847_n N_A_855_368#_M1003_g 0.0151225f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_733 N_A_1034_74#_c_837_n N_A_855_368#_M1003_g 0.00774077f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_734 N_A_1034_74#_c_860_n N_A_855_368#_M1003_g 0.00196389f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_735 N_A_1034_74#_c_847_n N_A_855_368#_c_1293_n 0.00483103f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_736 N_A_1034_74#_c_837_n N_A_855_368#_c_1293_n 0.0123734f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_737 N_A_1034_74#_c_850_n N_A_855_368#_c_1293_n 0.00422095f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_738 N_A_1034_74#_c_841_n N_A_855_368#_c_1293_n 0.00922521f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_739 N_A_1034_74#_c_826_n N_A_855_368#_c_1294_n 0.00922521f $X=9.085 $Y=1.16
+ $X2=0 $Y2=0
cc_740 N_A_1034_74#_c_842_n N_A_855_368#_c_1294_n 0.00132052f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_741 N_A_1034_74#_c_834_n N_A_855_368#_M1034_g 0.0039082f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_742 N_A_1034_74#_c_836_n N_A_855_368#_M1034_g 0.00172497f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_743 N_A_1034_74#_c_837_n N_A_855_368#_M1034_g 0.00175577f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_744 N_A_1034_74#_c_841_n N_A_855_368#_M1034_g 0.0213739f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_745 N_A_1034_74#_c_842_n N_A_855_368#_M1034_g 3.81838e-19 $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_746 N_A_1034_74#_c_829_n N_A_855_368#_c_1296_n 0.00513717f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_747 N_A_1034_74#_c_830_n N_A_855_368#_c_1296_n 0.00368996f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_748 N_A_1034_74#_c_839_n N_A_855_368#_c_1315_n 0.00764513f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_749 N_A_1034_74#_c_829_n N_A_855_368#_c_1298_n 0.00491662f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_750 N_A_1034_74#_c_829_n N_A_855_368#_c_1299_n 3.49166e-19 $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_751 N_A_1034_74#_c_839_n N_A_855_368#_c_1299_n 0.0122423f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_752 N_A_1034_74#_c_839_n N_A_855_368#_c_1317_n 0.00452944f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_753 N_A_1034_74#_c_829_n N_A_855_368#_c_1300_n 0.025108f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_754 N_A_1034_74#_c_838_n N_A_855_368#_c_1300_n 0.00839942f $X=5.382 $Y=1.075
+ $X2=0 $Y2=0
cc_755 N_A_1034_74#_c_839_n N_A_855_368#_c_1300_n 0.00962435f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_756 N_A_1034_74#_c_847_n N_A_2003_48#_c_1485_n 0.0213667f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_757 N_A_1034_74#_c_850_n N_A_2003_48#_c_1485_n 3.86848e-19 $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_758 N_A_1034_74#_c_847_n N_A_2003_48#_c_1494_n 0.0337241f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_759 N_A_1034_74#_c_834_n N_A_1745_74#_M1008_d 0.00191611f $X=8.825 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_760 N_A_1034_74#_c_836_n N_A_1745_74#_M1008_d 0.0113939f $X=8.91 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_761 N_A_1034_74#_c_842_n N_A_1745_74#_M1008_d 0.00132295f $X=9.33 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_762 N_A_1034_74#_c_837_n N_A_1745_74#_M1003_d 0.00800505f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_763 N_A_1034_74#_c_860_n N_A_1745_74#_M1003_d 0.00493868f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_764 N_A_1034_74#_c_850_n N_A_1745_74#_M1003_d 0.0018712f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_765 N_A_1034_74#_c_825_n N_A_1745_74#_c_1626_n 6.35408e-19 $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_766 N_A_1034_74#_c_834_n N_A_1745_74#_c_1626_n 0.00169523f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_767 N_A_1034_74#_c_836_n N_A_1745_74#_c_1626_n 0.0248143f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_768 N_A_1034_74#_c_841_n N_A_1745_74#_c_1626_n 0.00569557f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_769 N_A_1034_74#_c_842_n N_A_1745_74#_c_1626_n 0.0194065f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_770 N_A_1034_74#_c_847_n N_A_1745_74#_c_1595_n 0.0210277f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_771 N_A_1034_74#_c_860_n N_A_1745_74#_c_1595_n 0.0118084f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_772 N_A_1034_74#_c_850_n N_A_1745_74#_c_1595_n 0.0365613f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_773 N_A_1034_74#_c_836_n N_A_1745_74#_c_1582_n 0.00376918f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_774 N_A_1034_74#_c_837_n N_A_1745_74#_c_1583_n 0.0357282f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_775 N_A_1034_74#_c_841_n N_A_1745_74#_c_1583_n 5.18898e-19 $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_776 N_A_1034_74#_c_842_n N_A_1745_74#_c_1583_n 0.014106f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_777 N_A_1034_74#_c_847_n N_A_1745_74#_c_1597_n 0.00349139f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_778 N_A_1034_74#_c_850_n N_A_1745_74#_c_1597_n 0.0123723f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_779 N_A_1034_74#_c_847_n N_A_1745_74#_c_1598_n 9.40099e-19 $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_780 N_A_1034_74#_c_837_n N_A_1745_74#_c_1598_n 0.0141964f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_781 N_A_1034_74#_c_850_n N_A_1745_74#_c_1598_n 0.0119213f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_782 N_A_1034_74#_c_847_n N_A_1745_74#_c_1599_n 0.00429238f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_783 N_A_1034_74#_c_850_n N_A_1745_74#_c_1599_n 0.0246458f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_784 N_A_1034_74#_c_836_n N_A_1745_74#_c_1585_n 7.09256e-19 $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_785 N_A_1034_74#_c_841_n N_A_1745_74#_c_1585_n 5.62433e-19 $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_786 N_A_1034_74#_c_842_n N_A_1745_74#_c_1585_n 0.0131492f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_787 N_A_1034_74#_c_847_n N_VPWR_c_1869_n 0.00304676f $X=9.835 $Y=2.465 $X2=0
+ $Y2=0
cc_788 N_A_1034_74#_c_845_n N_VPWR_c_1854_n 9.39239e-19 $X=6.135 $Y=2.24 $X2=0
+ $Y2=0
cc_789 N_A_1034_74#_c_847_n N_VPWR_c_1854_n 0.00375679f $X=9.835 $Y=2.465 $X2=0
+ $Y2=0
cc_790 N_A_1034_74#_M1031_d N_A_415_81#_c_2053_n 0.00696197f $X=5.17 $Y=1.84
+ $X2=0 $Y2=0
cc_791 N_A_1034_74#_c_832_n N_A_415_81#_c_2053_n 0.00197233f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_792 N_A_1034_74#_c_839_n N_A_415_81#_c_2053_n 0.0224331f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_793 N_A_1034_74#_M1016_g N_A_415_81#_c_2047_n 2.10665e-19 $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_794 N_A_1034_74#_c_828_n N_A_415_81#_c_2047_n 0.0448129f $X=5.31 $Y=0.515
+ $X2=0 $Y2=0
cc_795 N_A_1034_74#_c_830_n N_A_415_81#_c_2047_n 0.0134743f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_796 N_A_1034_74#_M1016_g N_A_415_81#_c_2048_n 0.00683153f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_797 N_A_1034_74#_c_832_n N_A_415_81#_c_2048_n 0.0178348f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_798 N_A_1034_74#_c_843_n N_A_415_81#_c_2048_n 0.00650808f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_799 N_A_1034_74#_c_829_n N_A_415_81#_c_2049_n 0.0132327f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_800 N_A_1034_74#_c_832_n N_A_415_81#_c_2049_n 0.0143284f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_801 N_A_1034_74#_c_843_n N_A_415_81#_c_2049_n 3.9199e-19 $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_802 N_A_1034_74#_c_844_n N_A_415_81#_c_2055_n 0.00347407f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_803 N_A_1034_74#_c_845_n N_A_415_81#_c_2055_n 0.0091232f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_804 N_A_1034_74#_c_823_n N_A_415_81#_c_2055_n 0.00252722f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_805 N_A_1034_74#_c_832_n N_A_415_81#_c_2055_n 0.00801159f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_806 N_A_1034_74#_c_844_n N_A_415_81#_c_2050_n 0.00366894f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_807 N_A_1034_74#_c_823_n N_A_415_81#_c_2050_n 0.0104145f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_808 N_A_1034_74#_M1016_g N_A_415_81#_c_2050_n 0.00514657f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_809 N_A_1034_74#_c_832_n N_A_415_81#_c_2050_n 0.0256546f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_810 N_A_1034_74#_c_843_n N_A_415_81#_c_2050_n 0.00187233f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_811 N_A_1034_74#_c_844_n N_A_415_81#_c_2058_n 0.00129962f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_812 N_A_1034_74#_c_845_n N_A_415_81#_c_2058_n 0.0100992f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_813 N_A_1034_74#_c_832_n N_A_415_81#_c_2058_n 0.0221691f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_814 N_A_1034_74#_c_839_n N_A_415_81#_c_2058_n 0.00808762f $X=5.387 $Y=1.75
+ $X2=0 $Y2=0
cc_815 N_A_1034_74#_c_843_n N_A_415_81#_c_2058_n 0.00323194f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_816 N_A_1034_74#_c_833_n N_VGND_M1030_d 0.0162233f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_817 N_A_1034_74#_c_858_n N_VGND_M1030_d 0.00541973f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_818 N_A_1034_74#_c_835_n N_VGND_M1030_d 0.0011204f $X=8.1 $Y=0.34 $X2=0 $Y2=0
cc_819 N_A_1034_74#_c_831_n N_VGND_c_2262_n 0.00833854f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_820 N_A_1034_74#_c_830_n N_VGND_c_2272_n 0.0628549f $X=7.055 $Y=0.415 $X2=0
+ $Y2=0
cc_821 N_A_1034_74#_c_831_n N_VGND_c_2272_n 0.0229629f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_822 N_A_1034_74#_c_833_n N_VGND_c_2272_n 0.00392706f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_823 N_A_1034_74#_c_840_n N_VGND_c_2272_n 0.00787014f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_824 N_A_1034_74#_c_825_n N_VGND_c_2273_n 0.00278271f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_825 N_A_1034_74#_c_833_n N_VGND_c_2273_n 0.00335833f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_826 N_A_1034_74#_c_834_n N_VGND_c_2273_n 0.0579202f $X=8.825 $Y=0.34 $X2=0
+ $Y2=0
cc_827 N_A_1034_74#_c_835_n N_VGND_c_2273_n 0.0118998f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_828 N_A_1034_74#_c_833_n N_VGND_c_2277_n 0.0246013f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_829 N_A_1034_74#_c_835_n N_VGND_c_2277_n 0.0135791f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_830 N_A_1034_74#_c_840_n N_VGND_c_2277_n 0.00556242f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_831 N_A_1034_74#_c_825_n N_VGND_c_2282_n 0.00358928f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_832 N_A_1034_74#_c_830_n N_VGND_c_2282_n 0.0514347f $X=7.055 $Y=0.415 $X2=0
+ $Y2=0
cc_833 N_A_1034_74#_c_831_n N_VGND_c_2282_n 0.017632f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_834 N_A_1034_74#_c_833_n N_VGND_c_2282_n 0.0127392f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_835 N_A_1034_74#_c_834_n N_VGND_c_2282_n 0.0324872f $X=8.825 $Y=0.34 $X2=0
+ $Y2=0
cc_836 N_A_1034_74#_c_835_n N_VGND_c_2282_n 0.00655543f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_837 N_A_1034_74#_c_840_n N_VGND_c_2282_n 0.00618366f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_838 N_A_1034_74#_c_840_n A_1397_138# 0.00203667f $X=7.14 $Y=0.415 $X2=-0.19
+ $Y2=-0.245
cc_839 N_A_1367_112#_c_1046_n N_A_1233_138#_M1025_g 0.00313626f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_840 N_A_1367_112#_c_1070_n N_A_1233_138#_M1025_g 0.0131882f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_841 N_A_1367_112#_c_1046_n N_A_1233_138#_c_1153_n 0.00107505f $X=8.57
+ $Y=1.405 $X2=0 $Y2=0
cc_842 N_A_1367_112#_c_1047_n N_A_1233_138#_c_1153_n 0.0131822f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_843 N_A_1367_112#_c_1053_n N_A_1233_138#_c_1153_n 0.00530481f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_844 N_A_1367_112#_c_1094_n N_A_1233_138#_c_1153_n 0.00405015f $X=8.57
+ $Y=0.842 $X2=0 $Y2=0
cc_845 N_A_1367_112#_c_1053_n N_A_1233_138#_c_1161_n 0.0151257f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_846 N_A_1367_112#_M1001_g N_A_1233_138#_c_1171_n 0.004781f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_847 N_A_1367_112#_c_1067_n N_A_1233_138#_c_1171_n 0.0130756f $X=7.325
+ $Y=1.005 $X2=0 $Y2=0
cc_848 N_A_1367_112#_M1001_g N_A_1233_138#_c_1154_n 0.0095753f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_849 N_A_1367_112#_c_1048_n N_A_1233_138#_c_1154_n 0.0045184f $X=7.025 $Y=2.15
+ $X2=0 $Y2=0
cc_850 N_A_1367_112#_c_1049_n N_A_1233_138#_c_1154_n 9.21498e-19 $X=7.025
+ $Y=2.24 $X2=0 $Y2=0
cc_851 N_A_1367_112#_c_1044_n N_A_1233_138#_c_1154_n 0.062072f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_852 N_A_1367_112#_c_1045_n N_A_1233_138#_c_1154_n 0.0104616f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_853 N_A_1367_112#_c_1067_n N_A_1233_138#_c_1154_n 0.00114989f $X=7.325
+ $Y=1.005 $X2=0 $Y2=0
cc_854 N_A_1367_112#_c_1049_n N_A_1233_138#_c_1174_n 0.0109144f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_855 N_A_1367_112#_c_1044_n N_A_1233_138#_c_1174_n 0.00526266f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_856 N_A_1367_112#_c_1045_n N_A_1233_138#_c_1174_n 0.00311782f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_857 N_A_1367_112#_c_1048_n N_A_1233_138#_c_1155_n 0.00204704f $X=7.025
+ $Y=2.15 $X2=0 $Y2=0
cc_858 N_A_1367_112#_c_1049_n N_A_1233_138#_c_1155_n 0.00139157f $X=7.025
+ $Y=2.24 $X2=0 $Y2=0
cc_859 N_A_1367_112#_c_1044_n N_A_1233_138#_c_1155_n 0.0274325f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_860 N_A_1367_112#_c_1045_n N_A_1233_138#_c_1155_n 0.00208168f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_861 N_A_1367_112#_c_1044_n N_A_1233_138#_c_1156_n 0.0268297f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_862 N_A_1367_112#_c_1070_n N_A_1233_138#_c_1156_n 0.0133196f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_863 N_A_1367_112#_c_1046_n N_A_1233_138#_c_1157_n 0.0115079f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_864 N_A_1367_112#_c_1047_n N_A_1233_138#_c_1157_n 0.0142233f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_865 N_A_1367_112#_c_1070_n N_A_1233_138#_c_1157_n 0.0443118f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_866 N_A_1367_112#_c_1046_n N_A_1233_138#_c_1158_n 0.00161618f $X=8.57
+ $Y=1.405 $X2=0 $Y2=0
cc_867 N_A_1367_112#_c_1047_n N_A_1233_138#_c_1158_n 3.02987e-19 $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_868 N_A_1367_112#_c_1070_n N_A_1233_138#_c_1158_n 0.00252719f $X=8.27
+ $Y=0.842 $X2=0 $Y2=0
cc_869 N_A_1367_112#_c_1094_n N_A_1233_138#_c_1158_n 0.00137742f $X=8.57
+ $Y=0.842 $X2=0 $Y2=0
cc_870 N_A_1367_112#_M1001_g N_A_1233_138#_c_1159_n 0.00108413f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_871 N_A_1367_112#_c_1049_n N_A_1233_138#_c_1166_n 0.0060004f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_872 N_A_1367_112#_c_1049_n N_A_855_368#_c_1305_n 0.00323347f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_873 N_A_1367_112#_c_1049_n N_A_855_368#_c_1307_n 0.0307207f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_874 N_A_1367_112#_c_1049_n N_A_855_368#_c_1308_n 0.0100502f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_875 N_A_1367_112#_c_1053_n N_A_855_368#_c_1308_n 0.00400096f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_876 N_A_1367_112#_c_1053_n N_A_855_368#_c_1309_n 5.08057e-19 $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_877 N_A_1367_112#_c_1053_n N_A_855_368#_M1003_g 0.014001f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_878 N_A_1367_112#_c_1047_n N_A_855_368#_c_1294_n 0.0021457f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_879 N_A_1367_112#_c_1053_n N_A_855_368#_c_1294_n 0.00289869f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_880 N_A_1367_112#_c_1053_n N_A_1745_74#_c_1595_n 0.0146147f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_881 N_A_1367_112#_c_1049_n N_VPWR_c_1857_n 0.00433246f $X=7.025 $Y=2.24 $X2=0
+ $Y2=0
cc_882 N_A_1367_112#_c_1047_n N_VPWR_c_1859_n 0.00369686f $X=8.9 $Y=1.575 $X2=0
+ $Y2=0
cc_883 N_A_1367_112#_c_1053_n N_VPWR_c_1859_n 0.064586f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_884 N_A_1367_112#_c_1094_n N_VPWR_c_1859_n 0.00374786f $X=8.57 $Y=0.842 $X2=0
+ $Y2=0
cc_885 N_A_1367_112#_c_1053_n N_VPWR_c_1869_n 0.00748753f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_886 N_A_1367_112#_c_1049_n N_VPWR_c_1854_n 9.39239e-19 $X=7.025 $Y=2.24 $X2=0
+ $Y2=0
cc_887 N_A_1367_112#_c_1053_n N_VPWR_c_1854_n 0.00904755f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_888 N_A_1367_112#_M1001_g N_A_415_81#_c_2050_n 3.0177e-19 $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_889 N_A_1367_112#_c_1045_n N_A_415_81#_c_2050_n 6.15582e-19 $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_890 N_A_1367_112#_c_1070_n N_VGND_M1030_d 0.0155117f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_891 N_A_1367_112#_c_1067_n A_1397_138# 0.00267137f $X=7.325 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_892 N_A_1233_138#_c_1162_n N_A_855_368#_c_1303_n 0.00405916f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_893 N_A_1233_138#_c_1159_n N_A_855_368#_c_1292_n 0.00526454f $X=6.305 $Y=0.87
+ $X2=0 $Y2=0
cc_894 N_A_1233_138#_c_1162_n N_A_855_368#_c_1305_n 6.3693e-19 $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_895 N_A_1233_138#_c_1166_n N_A_855_368#_c_1305_n 3.29021e-19 $X=6.8 $Y=2.537
+ $X2=0 $Y2=0
cc_896 N_A_1233_138#_c_1162_n N_A_855_368#_c_1307_n 0.0128095f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_897 N_A_1233_138#_c_1154_n N_A_855_368#_c_1307_n 0.00130784f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_898 N_A_1233_138#_c_1161_n N_A_855_368#_c_1308_n 0.0103487f $X=8.675 $Y=1.66
+ $X2=0 $Y2=0
cc_899 N_A_1233_138#_c_1174_n N_A_855_368#_c_1308_n 0.00319775f $X=7.495
+ $Y=2.405 $X2=0 $Y2=0
cc_900 N_A_1233_138#_c_1155_n N_A_855_368#_c_1308_n 0.00775183f $X=7.58 $Y=2.32
+ $X2=0 $Y2=0
cc_901 N_A_1233_138#_c_1166_n N_A_855_368#_c_1308_n 0.00142193f $X=6.8 $Y=2.537
+ $X2=0 $Y2=0
cc_902 N_A_1233_138#_c_1161_n N_A_855_368#_c_1309_n 0.00230914f $X=8.675 $Y=1.66
+ $X2=0 $Y2=0
cc_903 N_A_1233_138#_c_1161_n N_A_855_368#_M1003_g 0.00599467f $X=8.675 $Y=1.66
+ $X2=0 $Y2=0
cc_904 N_A_1233_138#_c_1153_n N_A_855_368#_c_1294_n 0.00718094f $X=8.585 $Y=1.52
+ $X2=0 $Y2=0
cc_905 N_A_1233_138#_c_1174_n N_VPWR_M1032_d 0.00824542f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_906 N_A_1233_138#_c_1155_n N_VPWR_M1032_d 3.72881e-19 $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_907 N_A_1233_138#_c_1174_n N_VPWR_c_1857_n 0.0249179f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_908 N_A_1233_138#_c_1155_n N_VPWR_c_1857_n 0.00848094f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_909 N_A_1233_138#_c_1166_n N_VPWR_c_1857_n 0.00558555f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_910 N_A_1233_138#_c_1155_n N_VPWR_c_1858_n 0.00731736f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_911 N_A_1233_138#_c_1153_n N_VPWR_c_1859_n 0.00426403f $X=8.585 $Y=1.52 $X2=0
+ $Y2=0
cc_912 N_A_1233_138#_c_1161_n N_VPWR_c_1859_n 0.00771875f $X=8.675 $Y=1.66 $X2=0
+ $Y2=0
cc_913 N_A_1233_138#_c_1155_n N_VPWR_c_1859_n 0.0227303f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_914 N_A_1233_138#_c_1162_n N_VPWR_c_1873_n 0.00990874f $X=6.715 $Y=2.59 $X2=0
+ $Y2=0
cc_915 N_A_1233_138#_c_1166_n N_VPWR_c_1873_n 0.00390498f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_916 N_A_1233_138#_c_1161_n N_VPWR_c_1854_n 9.39239e-19 $X=8.675 $Y=1.66 $X2=0
+ $Y2=0
cc_917 N_A_1233_138#_c_1162_n N_VPWR_c_1854_n 0.0123809f $X=6.715 $Y=2.59 $X2=0
+ $Y2=0
cc_918 N_A_1233_138#_c_1174_n N_VPWR_c_1854_n 0.00931484f $X=7.495 $Y=2.405
+ $X2=0 $Y2=0
cc_919 N_A_1233_138#_c_1155_n N_VPWR_c_1854_n 0.0155791f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_920 N_A_1233_138#_c_1166_n N_VPWR_c_1854_n 0.00468883f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_921 N_A_1233_138#_c_1159_n N_A_415_81#_c_2047_n 0.0152023f $X=6.305 $Y=0.87
+ $X2=0 $Y2=0
cc_922 N_A_1233_138#_c_1171_n N_A_415_81#_c_2048_n 0.00571315f $X=6.715 $Y=0.99
+ $X2=0 $Y2=0
cc_923 N_A_1233_138#_c_1154_n N_A_415_81#_c_2048_n 0.0135849f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_924 N_A_1233_138#_c_1159_n N_A_415_81#_c_2048_n 0.021789f $X=6.305 $Y=0.87
+ $X2=0 $Y2=0
cc_925 N_A_1233_138#_c_1162_n N_A_415_81#_c_2055_n 0.0210559f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_926 N_A_1233_138#_c_1154_n N_A_415_81#_c_2055_n 0.0137319f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_927 N_A_1233_138#_c_1154_n N_A_415_81#_c_2050_n 0.048566f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_928 N_A_1233_138#_c_1162_n N_A_415_81#_c_2058_n 0.0131973f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_929 N_A_1233_138#_c_1154_n N_A_415_81#_c_2058_n 0.00169017f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_930 N_A_1233_138#_c_1166_n A_1342_463# 0.00298041f $X=6.8 $Y=2.537 $X2=-0.19
+ $Y2=-0.245
cc_931 N_A_1233_138#_M1025_g N_VGND_c_2273_n 0.00278271f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_932 N_A_1233_138#_M1025_g N_VGND_c_2277_n 0.00118431f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_933 N_A_1233_138#_M1025_g N_VGND_c_2282_n 0.00358928f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_934 N_A_1233_138#_c_1171_n A_1319_138# 0.00443085f $X=6.715 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_935 N_A_1233_138#_c_1154_n A_1319_138# 3.82916e-19 $X=6.8 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_936 N_A_855_368#_M1034_g N_A_2003_48#_M1028_g 0.0336121f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_937 N_A_855_368#_c_1293_n N_A_2003_48#_c_1485_n 0.00387806f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_938 N_A_855_368#_M1034_g N_A_2003_48#_c_1489_n 0.00111235f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_939 N_A_855_368#_c_1293_n N_A_2003_48#_c_1490_n 0.0336121f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_940 N_A_855_368#_M1034_g N_A_1745_74#_c_1626_n 0.0163048f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_941 N_A_855_368#_c_1309_n N_A_1745_74#_c_1595_n 0.00242116f $X=9.125 $Y=2.9
+ $X2=0 $Y2=0
cc_942 N_A_855_368#_M1003_g N_A_1745_74#_c_1595_n 0.00427038f $X=9.125 $Y=2.235
+ $X2=0 $Y2=0
cc_943 N_A_855_368#_M1034_g N_A_1745_74#_c_1582_n 0.00585097f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_944 N_A_855_368#_c_1293_n N_A_1745_74#_c_1583_n 0.00934901f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_945 N_A_855_368#_M1034_g N_A_1745_74#_c_1583_n 0.0140808f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_946 N_A_855_368#_M1034_g N_A_1745_74#_c_1584_n 0.00333053f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_947 N_A_855_368#_c_1293_n N_A_1745_74#_c_1597_n 3.21304e-19 $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_948 N_A_855_368#_M1034_g N_A_1745_74#_c_1585_n 0.00274755f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_949 N_A_855_368#_c_1315_n N_VPWR_M1019_d 0.0023273f $X=4.805 $Y=1.905 $X2=0
+ $Y2=0
cc_950 N_A_855_368#_c_1288_n N_VPWR_c_1856_n 0.00888208f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_951 N_A_855_368#_c_1290_n N_VPWR_c_1856_n 0.0017658f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_952 N_A_855_368#_c_1304_n N_VPWR_c_1856_n 0.00232909f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_953 N_A_855_368#_c_1305_n N_VPWR_c_1857_n 0.0060536f $X=6.635 $Y=2.9 $X2=0
+ $Y2=0
cc_954 N_A_855_368#_c_1308_n N_VPWR_c_1857_n 0.0264476f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_955 N_A_855_368#_c_1308_n N_VPWR_c_1858_n 0.0260616f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_956 N_A_855_368#_c_1308_n N_VPWR_c_1859_n 0.0170937f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_957 N_A_855_368#_c_1309_n N_VPWR_c_1859_n 0.00527525f $X=9.125 $Y=2.9 $X2=0
+ $Y2=0
cc_958 N_A_855_368#_c_1308_n N_VPWR_c_1869_n 0.0212209f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_959 N_A_855_368#_c_1288_n N_VPWR_c_1873_n 0.00413917f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_960 N_A_855_368#_c_1304_n N_VPWR_c_1873_n 0.0487125f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_961 N_A_855_368#_c_1288_n N_VPWR_c_1854_n 0.00399275f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_962 N_A_855_368#_c_1303_n N_VPWR_c_1854_n 0.024517f $X=6.545 $Y=3.15 $X2=0
+ $Y2=0
cc_963 N_A_855_368#_c_1304_n N_VPWR_c_1854_n 0.00693725f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_964 N_A_855_368#_c_1308_n N_VPWR_c_1854_n 0.0714547f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_965 N_A_855_368#_c_1314_n N_VPWR_c_1854_n 0.00495681f $X=6.635 $Y=3.15 $X2=0
+ $Y2=0
cc_966 N_A_855_368#_M1019_s N_A_415_81#_c_2053_n 0.0082239f $X=4.275 $Y=1.84
+ $X2=0 $Y2=0
cc_967 N_A_855_368#_c_1288_n N_A_415_81#_c_2053_n 0.0125758f $X=5.095 $Y=1.765
+ $X2=0 $Y2=0
cc_968 N_A_855_368#_c_1290_n N_A_415_81#_c_2053_n 0.0126563f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_969 N_A_855_368#_c_1315_n N_A_415_81#_c_2053_n 0.00790211f $X=4.805 $Y=1.905
+ $X2=0 $Y2=0
cc_970 N_A_855_368#_c_1317_n N_A_415_81#_c_2053_n 0.013838f $X=4.46 $Y=1.905
+ $X2=0 $Y2=0
cc_971 N_A_855_368#_c_1287_n N_A_415_81#_c_2047_n 4.04646e-19 $X=5.095 $Y=1.195
+ $X2=0 $Y2=0
cc_972 N_A_855_368#_c_1291_n N_A_415_81#_c_2047_n 0.0052952f $X=6.015 $Y=1.27
+ $X2=0 $Y2=0
cc_973 N_A_855_368#_c_1292_n N_A_415_81#_c_2047_n 0.00427356f $X=6.09 $Y=1.195
+ $X2=0 $Y2=0
cc_974 N_A_855_368#_c_1291_n N_A_415_81#_c_2048_n 0.0121754f $X=6.015 $Y=1.27
+ $X2=0 $Y2=0
cc_975 N_A_855_368#_c_1291_n N_A_415_81#_c_2049_n 0.00499805f $X=6.015 $Y=1.27
+ $X2=0 $Y2=0
cc_976 N_A_855_368#_c_1307_n N_A_415_81#_c_2055_n 6.45394e-19 $X=6.635 $Y=2.81
+ $X2=0 $Y2=0
cc_977 N_A_855_368#_c_1290_n N_A_415_81#_c_2050_n 0.00307189f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_978 N_A_855_368#_c_1290_n N_A_415_81#_c_2058_n 0.01209f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_979 N_A_855_368#_c_1303_n N_A_415_81#_c_2058_n 0.00570072f $X=6.545 $Y=3.15
+ $X2=0 $Y2=0
cc_980 N_A_855_368#_c_1307_n N_A_415_81#_c_2058_n 5.36672e-19 $X=6.635 $Y=2.81
+ $X2=0 $Y2=0
cc_981 N_A_855_368#_c_1339_n N_VGND_M1007_d 0.00226632f $X=4.805 $Y=1.005 $X2=0
+ $Y2=0
cc_982 N_A_855_368#_c_1298_n N_VGND_M1007_d 2.09292e-19 $X=4.89 $Y=1.245 $X2=0
+ $Y2=0
cc_983 N_A_855_368#_c_1297_n N_VGND_c_2261_n 0.0203528f $X=4.45 $Y=0.515 $X2=0
+ $Y2=0
cc_984 N_A_855_368#_c_1287_n N_VGND_c_2262_n 0.00260307f $X=5.095 $Y=1.195 $X2=0
+ $Y2=0
cc_985 N_A_855_368#_c_1297_n N_VGND_c_2262_n 0.0144259f $X=4.45 $Y=0.515 $X2=0
+ $Y2=0
cc_986 N_A_855_368#_c_1339_n N_VGND_c_2262_n 0.0159541f $X=4.805 $Y=1.005 $X2=0
+ $Y2=0
cc_987 N_A_855_368#_M1034_g N_VGND_c_2263_n 0.00156589f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_988 N_A_855_368#_c_1297_n N_VGND_c_2269_n 0.00749631f $X=4.45 $Y=0.515 $X2=0
+ $Y2=0
cc_989 N_A_855_368#_c_1287_n N_VGND_c_2272_n 0.00432683f $X=5.095 $Y=1.195 $X2=0
+ $Y2=0
cc_990 N_A_855_368#_M1034_g N_VGND_c_2273_n 0.00320499f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_991 N_A_855_368#_c_1287_n N_VGND_c_2282_n 0.00821393f $X=5.095 $Y=1.195 $X2=0
+ $Y2=0
cc_992 N_A_855_368#_M1034_g N_VGND_c_2282_n 0.00443186f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_993 N_A_855_368#_c_1297_n N_VGND_c_2282_n 0.0062048f $X=4.45 $Y=0.515 $X2=0
+ $Y2=0
cc_994 N_A_2003_48#_c_1487_n N_A_1745_74#_c_1573_n 0.00593167f $X=11.415 $Y=0.55
+ $X2=0 $Y2=0
cc_995 N_A_2003_48#_c_1488_n N_A_1745_74#_c_1573_n 0.00443992f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_996 N_A_2003_48#_c_1492_n N_A_1745_74#_c_1574_n 0.00146716f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_997 N_A_2003_48#_c_1491_n N_A_1745_74#_c_1590_n 0.00555199f $X=11.165 $Y=2.52
+ $X2=0 $Y2=0
cc_998 N_A_2003_48#_c_1488_n N_A_1745_74#_c_1575_n 0.00271488f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_999 N_A_2003_48#_c_1492_n N_A_1745_74#_c_1577_n 4.51356e-19 $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_1000 N_A_2003_48#_c_1488_n N_A_1745_74#_c_1579_n 0.00311356f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1001 N_A_2003_48#_c_1491_n N_A_1745_74#_c_1579_n 0.0136035f $X=11.165 $Y=2.52
+ $X2=0 $Y2=0
cc_1002 N_A_2003_48#_c_1492_n N_A_1745_74#_c_1579_n 0.0149058f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_1003 N_A_2003_48#_M1028_g N_A_1745_74#_c_1626_n 0.00125881f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_1004 N_A_2003_48#_c_1494_n N_A_1745_74#_c_1595_n 0.0108165f $X=10.255
+ $Y=2.465 $X2=0 $Y2=0
cc_1005 N_A_2003_48#_M1028_g N_A_1745_74#_c_1582_n 9.29499e-19 $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_1006 N_A_2003_48#_M1028_g N_A_1745_74#_c_1583_n 0.00223708f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_1007 N_A_2003_48#_c_1485_n N_A_1745_74#_c_1583_n 0.00234903f $X=10.255
+ $Y=2.375 $X2=0 $Y2=0
cc_1008 N_A_2003_48#_c_1489_n N_A_1745_74#_c_1583_n 0.0167585f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1009 N_A_2003_48#_M1028_g N_A_1745_74#_c_1584_n 0.0143799f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_1010 N_A_2003_48#_c_1486_n N_A_1745_74#_c_1584_n 0.0259611f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_1011 N_A_2003_48#_c_1489_n N_A_1745_74#_c_1584_n 0.0242156f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1012 N_A_2003_48#_c_1490_n N_A_1745_74#_c_1584_n 0.001245f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1013 N_A_2003_48#_c_1485_n N_A_1745_74#_c_1597_n 0.00995549f $X=10.255
+ $Y=2.375 $X2=0 $Y2=0
cc_1014 N_A_2003_48#_c_1489_n N_A_1745_74#_c_1597_n 0.0210104f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1015 N_A_2003_48#_c_1490_n N_A_1745_74#_c_1597_n 0.00106876f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1016 N_A_2003_48#_c_1485_n N_A_1745_74#_c_1599_n 0.0141267f $X=10.255
+ $Y=2.375 $X2=0 $Y2=0
cc_1017 N_A_2003_48#_c_1494_n N_A_1745_74#_c_1599_n 0.00550853f $X=10.255
+ $Y=2.465 $X2=0 $Y2=0
cc_1018 N_A_2003_48#_c_1486_n N_A_1745_74#_c_1586_n 0.0247317f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_1019 N_A_2003_48#_c_1487_n N_A_1745_74#_c_1586_n 0.014253f $X=11.415 $Y=0.55
+ $X2=0 $Y2=0
cc_1020 N_A_2003_48#_c_1488_n N_A_1745_74#_c_1586_n 0.0236842f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1021 N_A_2003_48#_c_1486_n N_A_1745_74#_c_1587_n 0.0121221f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_1022 N_A_2003_48#_c_1487_n N_A_1745_74#_c_1587_n 0.00619797f $X=11.415
+ $Y=0.55 $X2=0 $Y2=0
cc_1023 N_A_2003_48#_c_1488_n N_A_1745_74#_c_1587_n 0.0191241f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1024 N_A_2003_48#_c_1487_n N_A_2339_74#_c_1743_n 0.026931f $X=11.415 $Y=0.55
+ $X2=0 $Y2=0
cc_1025 N_A_2003_48#_c_1488_n N_A_2339_74#_c_1743_n 0.0405862f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1026 N_A_2003_48#_c_1488_n N_A_2339_74#_c_1745_n 0.00909743f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1027 N_A_2003_48#_c_1491_n N_A_2339_74#_c_1745_n 0.00195796f $X=11.165
+ $Y=2.52 $X2=0 $Y2=0
cc_1028 N_A_2003_48#_c_1492_n N_A_2339_74#_c_1745_n 0.0157384f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_1029 N_A_2003_48#_c_1494_n N_VPWR_c_1860_n 0.00888901f $X=10.255 $Y=2.465
+ $X2=0 $Y2=0
cc_1030 N_A_2003_48#_c_1495_n N_VPWR_c_1860_n 0.0309795f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1031 N_A_2003_48#_c_1491_n N_VPWR_c_1861_n 0.057723f $X=11.165 $Y=2.52 $X2=0
+ $Y2=0
cc_1032 N_A_2003_48#_c_1494_n N_VPWR_c_1869_n 0.00341164f $X=10.255 $Y=2.465
+ $X2=0 $Y2=0
cc_1033 N_A_2003_48#_c_1495_n N_VPWR_c_1874_n 0.0143991f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1034 N_A_2003_48#_c_1494_n N_VPWR_c_1854_n 0.00538309f $X=10.255 $Y=2.465
+ $X2=0 $Y2=0
cc_1035 N_A_2003_48#_c_1495_n N_VPWR_c_1854_n 0.0119711f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1036 N_A_2003_48#_M1028_g N_VGND_c_2263_n 0.00986387f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1037 N_A_2003_48#_c_1487_n N_VGND_c_2263_n 0.0104724f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1038 N_A_2003_48#_M1028_g N_VGND_c_2273_n 0.00383152f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1039 N_A_2003_48#_c_1487_n N_VGND_c_2274_n 0.0191719f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1040 N_A_2003_48#_M1028_g N_VGND_c_2282_n 0.0075725f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1041 N_A_2003_48#_c_1487_n N_VGND_c_2282_n 0.0192149f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1042 N_A_1745_74#_c_1576_n N_A_2339_74#_c_1737_n 0.00970941f $X=12.055
+ $Y=1.185 $X2=0 $Y2=0
cc_1043 N_A_1745_74#_c_1578_n N_A_2339_74#_c_1739_n 0.00924572f $X=12.415
+ $Y=1.69 $X2=0 $Y2=0
cc_1044 N_A_1745_74#_c_1581_n N_A_2339_74#_c_1739_n 0.00970941f $X=12.055
+ $Y=1.26 $X2=0 $Y2=0
cc_1045 N_A_1745_74#_c_1593_n N_A_2339_74#_c_1748_n 0.0130951f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1046 N_A_1745_74#_c_1573_n N_A_2339_74#_c_1743_n 5.54394e-19 $X=10.99 $Y=0.9
+ $X2=0 $Y2=0
cc_1047 N_A_1745_74#_c_1575_n N_A_2339_74#_c_1743_n 0.00765913f $X=11.98 $Y=1.26
+ $X2=0 $Y2=0
cc_1048 N_A_1745_74#_c_1576_n N_A_2339_74#_c_1743_n 0.0035045f $X=12.055
+ $Y=1.185 $X2=0 $Y2=0
cc_1049 N_A_1745_74#_c_1587_n N_A_2339_74#_c_1743_n 8.98164e-19 $X=11.535
+ $Y=1.117 $X2=0 $Y2=0
cc_1050 N_A_1745_74#_c_1574_n N_A_2339_74#_c_1744_n 0.00115484f $X=11.475
+ $Y=1.665 $X2=0 $Y2=0
cc_1051 N_A_1745_74#_c_1591_n N_A_2339_74#_c_1744_n 0.0135732f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1052 N_A_1745_74#_c_1577_n N_A_2339_74#_c_1744_n 6.63362e-19 $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1053 N_A_1745_74#_c_1578_n N_A_2339_74#_c_1744_n 0.0137178f $X=12.415 $Y=1.69
+ $X2=0 $Y2=0
cc_1054 N_A_1745_74#_c_1593_n N_A_2339_74#_c_1744_n 0.0135773f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1055 N_A_1745_74#_c_1580_n N_A_2339_74#_c_1744_n 0.00313656f $X=12.04 $Y=1.69
+ $X2=0 $Y2=0
cc_1056 N_A_1745_74#_c_1574_n N_A_2339_74#_c_1745_n 2.72834e-19 $X=11.475
+ $Y=1.665 $X2=0 $Y2=0
cc_1057 N_A_1745_74#_c_1575_n N_A_2339_74#_c_1745_n 0.00807224f $X=11.98 $Y=1.26
+ $X2=0 $Y2=0
cc_1058 N_A_1745_74#_c_1577_n N_A_2339_74#_c_1745_n 0.0179017f $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1059 N_A_1745_74#_c_1578_n N_A_2339_74#_c_1745_n 0.00885109f $X=12.415
+ $Y=1.69 $X2=0 $Y2=0
cc_1060 N_A_1745_74#_c_1579_n N_A_2339_74#_c_1745_n 0.00110135f $X=11.475
+ $Y=1.575 $X2=0 $Y2=0
cc_1061 N_A_1745_74#_c_1580_n N_A_2339_74#_c_1745_n 0.00144773f $X=12.04 $Y=1.69
+ $X2=0 $Y2=0
cc_1062 N_A_1745_74#_c_1581_n N_A_2339_74#_c_1745_n 0.00802343f $X=12.055
+ $Y=1.26 $X2=0 $Y2=0
cc_1063 N_A_1745_74#_c_1577_n N_A_2339_74#_c_1747_n 0.00212764f $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1064 N_A_1745_74#_c_1578_n N_A_2339_74#_c_1747_n 0.00620598f $X=12.415
+ $Y=1.69 $X2=0 $Y2=0
cc_1065 N_A_1745_74#_c_1595_n N_VPWR_c_1860_n 0.0271933f $X=10.125 $Y=2.715
+ $X2=0 $Y2=0
cc_1066 N_A_1745_74#_c_1599_n N_VPWR_c_1860_n 0.00221611f $X=10.21 $Y=2.55 $X2=0
+ $Y2=0
cc_1067 N_A_1745_74#_c_1589_n N_VPWR_c_1861_n 0.0068494f $X=11.475 $Y=2.375
+ $X2=0 $Y2=0
cc_1068 N_A_1745_74#_c_1590_n N_VPWR_c_1861_n 0.0116785f $X=11.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1069 N_A_1745_74#_c_1575_n N_VPWR_c_1861_n 0.00368592f $X=11.98 $Y=1.26 $X2=0
+ $Y2=0
cc_1070 N_A_1745_74#_c_1591_n N_VPWR_c_1861_n 0.00713044f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1071 N_A_1745_74#_c_1593_n N_VPWR_c_1862_n 0.0107123f $X=12.49 $Y=1.765 $X2=0
+ $Y2=0
cc_1072 N_A_1745_74#_c_1595_n N_VPWR_c_1869_n 0.0274709f $X=10.125 $Y=2.715
+ $X2=0 $Y2=0
cc_1073 N_A_1745_74#_c_1590_n N_VPWR_c_1874_n 0.00461464f $X=11.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1074 N_A_1745_74#_c_1591_n N_VPWR_c_1875_n 0.00393873f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1075 N_A_1745_74#_c_1593_n N_VPWR_c_1875_n 0.00393873f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1076 N_A_1745_74#_c_1590_n N_VPWR_c_1854_n 0.00990964f $X=11.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1077 N_A_1745_74#_c_1591_n N_VPWR_c_1854_n 0.00462577f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1078 N_A_1745_74#_c_1593_n N_VPWR_c_1854_n 0.00462577f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1079 N_A_1745_74#_c_1595_n N_VPWR_c_1854_n 0.0333279f $X=10.125 $Y=2.715
+ $X2=0 $Y2=0
cc_1080 N_A_1745_74#_c_1595_n A_1982_508# 0.00498821f $X=10.125 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1081 N_A_1745_74#_c_1573_n N_VGND_c_2263_n 0.00154514f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1082 N_A_1745_74#_c_1626_n N_VGND_c_2263_n 0.011455f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1083 N_A_1745_74#_c_1584_n N_VGND_c_2263_n 0.0267689f $X=10.915 $Y=0.97 $X2=0
+ $Y2=0
cc_1084 N_A_1745_74#_c_1576_n N_VGND_c_2264_n 0.0149682f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1085 N_A_1745_74#_c_1626_n N_VGND_c_2273_n 0.0190071f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1086 N_A_1745_74#_c_1573_n N_VGND_c_2274_n 0.00433941f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1087 N_A_1745_74#_c_1576_n N_VGND_c_2274_n 0.00383152f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1088 N_A_1745_74#_c_1573_n N_VGND_c_2282_n 0.00822721f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1089 N_A_1745_74#_c_1576_n N_VGND_c_2282_n 0.00762539f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1090 N_A_1745_74#_c_1626_n N_VGND_c_2282_n 0.0200126f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1091 N_A_2339_74#_c_1744_n N_VPWR_c_1861_n 0.059064f $X=12.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1092 N_A_2339_74#_c_1745_n N_VPWR_c_1861_n 0.0106252f $X=12.43 $Y=1.435 $X2=0
+ $Y2=0
cc_1093 N_A_2339_74#_c_1738_n N_VPWR_c_1862_n 9.84896e-19 $X=12.84 $Y=1.3 $X2=0
+ $Y2=0
cc_1094 N_A_2339_74#_c_1748_n N_VPWR_c_1862_n 0.0091433f $X=13.025 $Y=1.765
+ $X2=0 $Y2=0
cc_1095 N_A_2339_74#_c_1744_n N_VPWR_c_1862_n 0.0579567f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1096 N_A_2339_74#_c_1746_n N_VPWR_c_1862_n 0.0181117f $X=13.685 $Y=1.435
+ $X2=0 $Y2=0
cc_1097 N_A_2339_74#_c_1747_n N_VPWR_c_1862_n 0.00116289f $X=14.375 $Y=1.495
+ $X2=0 $Y2=0
cc_1098 N_A_2339_74#_c_1748_n N_VPWR_c_1863_n 0.00445602f $X=13.025 $Y=1.765
+ $X2=0 $Y2=0
cc_1099 N_A_2339_74#_c_1749_n N_VPWR_c_1863_n 0.00445602f $X=13.475 $Y=1.765
+ $X2=0 $Y2=0
cc_1100 N_A_2339_74#_c_1749_n N_VPWR_c_1864_n 0.00653972f $X=13.475 $Y=1.765
+ $X2=0 $Y2=0
cc_1101 N_A_2339_74#_c_1750_n N_VPWR_c_1864_n 0.0140029f $X=13.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1102 N_A_2339_74#_c_1751_n N_VPWR_c_1864_n 5.97443e-19 $X=14.375 $Y=1.765
+ $X2=0 $Y2=0
cc_1103 N_A_2339_74#_c_1751_n N_VPWR_c_1866_n 0.00671837f $X=14.375 $Y=1.765
+ $X2=0 $Y2=0
cc_1104 N_A_2339_74#_c_1744_n N_VPWR_c_1875_n 0.00664674f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1105 N_A_2339_74#_c_1750_n N_VPWR_c_1876_n 0.00413917f $X=13.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1106 N_A_2339_74#_c_1751_n N_VPWR_c_1876_n 0.00461464f $X=14.375 $Y=1.765
+ $X2=0 $Y2=0
cc_1107 N_A_2339_74#_c_1748_n N_VPWR_c_1854_n 0.00862391f $X=13.025 $Y=1.765
+ $X2=0 $Y2=0
cc_1108 N_A_2339_74#_c_1749_n N_VPWR_c_1854_n 0.00857589f $X=13.475 $Y=1.765
+ $X2=0 $Y2=0
cc_1109 N_A_2339_74#_c_1750_n N_VPWR_c_1854_n 0.00817726f $X=13.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1110 N_A_2339_74#_c_1751_n N_VPWR_c_1854_n 0.00911437f $X=14.375 $Y=1.765
+ $X2=0 $Y2=0
cc_1111 N_A_2339_74#_c_1744_n N_VPWR_c_1854_n 0.00995652f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1112 N_A_2339_74#_c_1737_n N_Q_c_2193_n 0.00667713f $X=12.485 $Y=1.225 $X2=0
+ $Y2=0
cc_1113 N_A_2339_74#_c_1740_n N_Q_c_2193_n 0.0125407f $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1114 N_A_2339_74#_c_1740_n N_Q_c_2204_n 0.0131906f $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1115 N_A_2339_74#_c_1741_n N_Q_c_2204_n 0.0164113f $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1116 N_A_2339_74#_c_1746_n N_Q_c_2204_n 0.0693421f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1117 N_A_2339_74#_c_1747_n N_Q_c_2204_n 0.0179128f $X=14.375 $Y=1.495 $X2=0
+ $Y2=0
cc_1118 N_A_2339_74#_c_1737_n N_Q_c_2208_n 0.00205797f $X=12.485 $Y=1.225 $X2=0
+ $Y2=0
cc_1119 N_A_2339_74#_c_1738_n N_Q_c_2208_n 0.00210982f $X=12.84 $Y=1.3 $X2=0
+ $Y2=0
cc_1120 N_A_2339_74#_c_1740_n N_Q_c_2208_n 7.32094e-19 $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1121 N_A_2339_74#_c_1746_n N_Q_c_2208_n 0.0218379f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1122 N_A_2339_74#_c_1748_n N_Q_c_2197_n 0.0117913f $X=13.025 $Y=1.765 $X2=0
+ $Y2=0
cc_1123 N_A_2339_74#_c_1749_n N_Q_c_2197_n 0.0130095f $X=13.475 $Y=1.765 $X2=0
+ $Y2=0
cc_1124 N_A_2339_74#_c_1750_n N_Q_c_2197_n 7.91051e-19 $X=13.925 $Y=1.765 $X2=0
+ $Y2=0
cc_1125 N_A_2339_74#_c_1749_n N_Q_c_2198_n 0.0120074f $X=13.475 $Y=1.765 $X2=0
+ $Y2=0
cc_1126 N_A_2339_74#_c_1750_n N_Q_c_2198_n 0.0157775f $X=13.925 $Y=1.765 $X2=0
+ $Y2=0
cc_1127 N_A_2339_74#_c_1746_n N_Q_c_2198_n 0.0321534f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1128 N_A_2339_74#_c_1747_n N_Q_c_2198_n 0.00943636f $X=14.375 $Y=1.495 $X2=0
+ $Y2=0
cc_1129 N_A_2339_74#_c_1748_n N_Q_c_2199_n 0.0033048f $X=13.025 $Y=1.765 $X2=0
+ $Y2=0
cc_1130 N_A_2339_74#_c_1749_n N_Q_c_2199_n 0.00132156f $X=13.475 $Y=1.765 $X2=0
+ $Y2=0
cc_1131 N_A_2339_74#_c_1744_n N_Q_c_2199_n 0.00129097f $X=12.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1132 N_A_2339_74#_c_1746_n N_Q_c_2199_n 0.0276943f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1133 N_A_2339_74#_c_1747_n N_Q_c_2199_n 0.00739484f $X=14.375 $Y=1.495 $X2=0
+ $Y2=0
cc_1134 N_A_2339_74#_c_1750_n N_Q_c_2200_n 0.00471332f $X=13.925 $Y=1.765 $X2=0
+ $Y2=0
cc_1135 N_A_2339_74#_c_1751_n N_Q_c_2200_n 4.03081e-19 $X=14.375 $Y=1.765 $X2=0
+ $Y2=0
cc_1136 N_A_2339_74#_c_1741_n N_Q_c_2194_n 3.92031e-19 $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1137 N_A_2339_74#_c_1742_n N_Q_c_2194_n 3.92313e-19 $X=14.385 $Y=1.225 $X2=0
+ $Y2=0
cc_1138 N_A_2339_74#_c_1741_n N_Q_c_2195_n 0.00272065f $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1139 N_A_2339_74#_c_1742_n N_Q_c_2195_n 0.00240279f $X=14.385 $Y=1.225 $X2=0
+ $Y2=0
cc_1140 N_A_2339_74#_c_1746_n N_Q_c_2195_n 0.00167694f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1141 N_A_2339_74#_c_1747_n N_Q_c_2195_n 0.00901833f $X=14.375 $Y=1.495 $X2=0
+ $Y2=0
cc_1142 N_A_2339_74#_c_1751_n Q 0.0145189f $X=14.375 $Y=1.765 $X2=0 $Y2=0
cc_1143 N_A_2339_74#_c_1746_n Q 0.0194661f $X=13.685 $Y=1.435 $X2=0 $Y2=0
cc_1144 N_A_2339_74#_c_1747_n Q 0.050284f $X=14.375 $Y=1.495 $X2=0 $Y2=0
cc_1145 N_A_2339_74#_c_1737_n N_VGND_c_2264_n 0.00182441f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1146 N_A_2339_74#_c_1743_n N_VGND_c_2264_n 0.0266033f $X=11.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1147 N_A_2339_74#_c_1745_n N_VGND_c_2264_n 0.0191073f $X=12.43 $Y=1.435 $X2=0
+ $Y2=0
cc_1148 N_A_2339_74#_c_1741_n N_VGND_c_2266_n 4.98647e-19 $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1149 N_A_2339_74#_c_1742_n N_VGND_c_2266_n 0.0149937f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1150 N_A_2339_74#_c_1743_n N_VGND_c_2274_n 0.00749631f $X=11.84 $Y=0.515
+ $X2=0 $Y2=0
cc_1151 N_A_2339_74#_c_1741_n N_VGND_c_2275_n 0.00383152f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1152 N_A_2339_74#_c_1742_n N_VGND_c_2275_n 0.00383152f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1153 N_A_2339_74#_c_1737_n N_VGND_c_2280_n 0.00434272f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1154 N_A_2339_74#_c_1740_n N_VGND_c_2280_n 0.00434272f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1155 N_A_2339_74#_c_1740_n N_VGND_c_2281_n 0.00452683f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1156 N_A_2339_74#_c_1741_n N_VGND_c_2281_n 0.0108787f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1157 N_A_2339_74#_c_1742_n N_VGND_c_2281_n 4.44374e-19 $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1158 N_A_2339_74#_c_1737_n N_VGND_c_2282_n 0.00820158f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1159 N_A_2339_74#_c_1740_n N_VGND_c_2282_n 0.00825037f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1160 N_A_2339_74#_c_1741_n N_VGND_c_2282_n 0.00752925f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1161 N_A_2339_74#_c_1742_n N_VGND_c_2282_n 0.0075754f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1162 N_A_2339_74#_c_1743_n N_VGND_c_2282_n 0.0062048f $X=11.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1163 N_VPWR_M1006_d N_A_415_81#_c_2059_n 0.0110267f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1164 N_VPWR_c_1855_n N_A_415_81#_c_2059_n 0.0214041f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1165 N_VPWR_c_1854_n N_A_415_81#_c_2059_n 0.0231955f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1166 N_VPWR_c_1855_n N_A_415_81#_c_2052_n 0.02127f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1167 N_VPWR_c_1867_n N_A_415_81#_c_2052_n 0.0166211f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1168 N_VPWR_c_1854_n N_A_415_81#_c_2052_n 0.0136307f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1169 N_VPWR_M1019_d N_A_415_81#_c_2053_n 0.00463341f $X=4.72 $Y=1.84 $X2=0
+ $Y2=0
cc_1170 N_VPWR_c_1856_n N_A_415_81#_c_2053_n 0.0166996f $X=4.87 $Y=2.815 $X2=0
+ $Y2=0
cc_1171 N_VPWR_c_1854_n N_A_415_81#_c_2053_n 0.0501229f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1172 N_VPWR_M1006_d N_A_415_81#_c_2054_n 8.56696e-19 $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1173 N_VPWR_c_1854_n N_A_415_81#_c_2054_n 0.00615626f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1174 N_VPWR_c_1855_n N_A_415_81#_c_2057_n 0.00713257f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1175 N_VPWR_c_1872_n N_A_415_81#_c_2057_n 0.0144799f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1176 N_VPWR_c_1877_n N_A_415_81#_c_2057_n 0.0198341f $X=1.4 $Y=2.465 $X2=0
+ $Y2=0
cc_1177 N_VPWR_c_1854_n N_A_415_81#_c_2057_n 0.0119509f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1178 N_VPWR_c_1873_n N_A_415_81#_c_2058_n 0.00751117f $X=7.17 $Y=3.33 $X2=0
+ $Y2=0
cc_1179 N_VPWR_c_1854_n N_A_415_81#_c_2058_n 0.00907713f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1180 N_VPWR_c_1862_n N_Q_c_2197_n 0.0697297f $X=12.8 $Y=1.985 $X2=0 $Y2=0
cc_1181 N_VPWR_c_1863_n N_Q_c_2197_n 0.014552f $X=13.615 $Y=3.33 $X2=0 $Y2=0
cc_1182 N_VPWR_c_1864_n N_Q_c_2197_n 0.058364f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1183 N_VPWR_c_1854_n N_Q_c_2197_n 0.0119791f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1184 N_VPWR_M1004_d N_Q_c_2198_n 0.00222494f $X=13.55 $Y=1.84 $X2=0 $Y2=0
cc_1185 N_VPWR_c_1864_n N_Q_c_2198_n 0.0154248f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1186 N_VPWR_c_1862_n N_Q_c_2199_n 0.00857239f $X=12.8 $Y=1.985 $X2=0 $Y2=0
cc_1187 N_VPWR_c_1864_n N_Q_c_2200_n 0.0565072f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1188 N_VPWR_c_1866_n N_Q_c_2200_n 0.00140347f $X=14.6 $Y=2.275 $X2=0 $Y2=0
cc_1189 N_VPWR_c_1876_n N_Q_c_2200_n 0.00950426f $X=14.47 $Y=3.33 $X2=0 $Y2=0
cc_1190 N_VPWR_c_1854_n N_Q_c_2200_n 0.0078668f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1191 N_VPWR_M1044_d Q 0.0031824f $X=14.45 $Y=1.84 $X2=0 $Y2=0
cc_1192 N_VPWR_c_1866_n Q 0.0222952f $X=14.6 $Y=2.275 $X2=0 $Y2=0
cc_1193 N_A_415_81#_c_2059_n A_514_464# 0.013941f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1194 N_A_415_81#_M1010_d N_noxref_24_c_2403_n 0.00945085f $X=2.075 $Y=0.405
+ $X2=0 $Y2=0
cc_1195 N_A_415_81#_c_2044_n N_noxref_24_c_2403_n 0.028856f $X=2.565 $Y=0.72
+ $X2=0 $Y2=0
cc_1196 N_A_415_81#_c_2045_n N_noxref_24_c_2403_n 0.0134817f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1197 N_A_415_81#_c_2044_n N_noxref_24_c_2405_n 0.00467283f $X=2.565 $Y=0.72
+ $X2=0 $Y2=0
cc_1198 N_A_415_81#_c_2045_n N_noxref_24_c_2405_n 0.0221136f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1199 N_Q_c_2204_n N_VGND_M1018_d 0.019527f $X=14.085 $Y=1.015 $X2=0 $Y2=0
cc_1200 N_Q_c_2193_n N_VGND_c_2264_n 0.0224879f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1201 N_Q_c_2194_n N_VGND_c_2266_n 0.0214745f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1202 N_Q_c_2195_n N_VGND_c_2266_n 0.00176181f $X=14.17 $Y=1.3 $X2=0 $Y2=0
cc_1203 Q N_VGND_c_2266_n 0.0295377f $X=14.555 $Y=1.58 $X2=0 $Y2=0
cc_1204 N_Q_c_2194_n N_VGND_c_2275_n 0.00749631f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1205 N_Q_c_2193_n N_VGND_c_2280_n 0.0144922f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1206 N_Q_c_2193_n N_VGND_c_2281_n 0.0163053f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1207 N_Q_c_2204_n N_VGND_c_2281_n 0.0647108f $X=14.085 $Y=1.015 $X2=0 $Y2=0
cc_1208 N_Q_c_2194_n N_VGND_c_2281_n 0.0171417f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1209 N_Q_c_2193_n N_VGND_c_2282_n 0.0118826f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1210 N_Q_c_2194_n N_VGND_c_2282_n 0.0062048f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1211 N_VGND_c_2267_n N_noxref_24_c_2403_n 0.115309f $X=3.725 $Y=0 $X2=0 $Y2=0
cc_1212 N_VGND_c_2282_n N_noxref_24_c_2403_n 0.0673001f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1213 N_VGND_c_2260_n N_noxref_24_c_2404_n 0.0259561f $X=0.71 $Y=0.555 $X2=0
+ $Y2=0
cc_1214 N_VGND_c_2267_n N_noxref_24_c_2404_n 0.0225398f $X=3.725 $Y=0 $X2=0
+ $Y2=0
cc_1215 N_VGND_c_2282_n N_noxref_24_c_2404_n 0.0125704f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1216 N_VGND_c_2261_n N_noxref_24_c_2405_n 0.0248556f $X=3.89 $Y=0.605 $X2=0
+ $Y2=0
cc_1217 N_VGND_c_2267_n N_noxref_24_c_2405_n 0.0229596f $X=3.725 $Y=0 $X2=0
+ $Y2=0
cc_1218 N_VGND_c_2282_n N_noxref_24_c_2405_n 0.0126481f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1219 N_noxref_24_c_2403_n noxref_25 0.00373495f $X=3.225 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1220 N_noxref_24_c_2403_n noxref_26 0.00226367f $X=3.225 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
