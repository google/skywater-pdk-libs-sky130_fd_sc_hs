* File: sky130_fd_sc_hs__nand3b_4.spice
* Created: Tue Sep  1 20:09:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nand3b_4.pex.spice"
.subckt sky130_fd_sc_hs__nand3b_4  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_N_M1000_g N_A_89_172#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.203425 AS=0.19515 PD=1.425 PS=2.05 NRD=35.652 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1004 N_A_297_82#_M1004_d N_C_M1004_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.203425 PD=1.02 PS=1.425 NRD=0 NRS=35.652 M=1 R=4.93333
+ SA=75000.8 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1009 N_A_297_82#_M1004_d N_C_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2715 PD=1.02 PS=1.56 NRD=0 NRS=50.568 M=1 R=4.93333 SA=75001.2
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1011 N_A_297_82#_M1011_d N_C_M1011_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2715 PD=1.09 PS=1.56 NRD=0 NRS=50.568 M=1 R=4.93333 SA=75002
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_A_297_82#_M1011_d N_C_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.19935 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_744_74#_M1002_d N_A_89_172#_M1002_g N_Y_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1962 AS=0.11285 PD=2.05 PS=1.045 NRD=0 NRS=1.62 M=1 R=4.93333
+ SA=75000.2 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1016 N_A_744_74#_M1016_d N_A_89_172#_M1016_g N_Y_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75000.6 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1017 N_A_744_74#_M1016_d N_A_89_172#_M1017_g N_Y_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1020 N_A_744_74#_M1020_d N_A_89_172#_M1020_g N_Y_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002 A=0.111 P=1.78 MULT=1
MM1001 N_A_744_74#_M1020_d N_B_M1001_g N_A_297_82#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1005 N_A_744_74#_M1005_d N_B_M1005_g N_A_297_82#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1018 N_A_744_74#_M1005_d N_B_M1018_g N_A_297_82#_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1019 N_A_744_74#_M1019_d N_B_M1019_g N_A_297_82#_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1976 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_89_172#_M1003_d N_A_N_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.5754 PD=1.14 PS=3.05 NRD=2.3443 NRS=93.7917 M=1 R=5.6 SA=75000.6
+ SB=75006.5 A=0.126 P=1.98 MULT=1
MM1006 N_A_89_172#_M1003_d N_A_N_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.5316 PD=1.14 PS=1.92857 NRD=2.3443 NRS=135.516 M=1 R=5.6
+ SA=75001.1 SB=75006 A=0.126 P=1.98 MULT=1
MM1010 N_Y_M1010_d N_C_M1010_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.7088 PD=1.42 PS=2.57143 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75004.8 A=0.168 P=2.54 MULT=1
MM1012 N_Y_M1010_d N_C_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.2604 PD=1.42 PS=1.585 NRD=1.7533 NRS=15.8191 M=1 R=7.46667 SA=75002.4
+ SB=75004.3 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1012_s N_A_89_172#_M1014_g N_Y_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2604 AS=0.3808 PD=1.585 PS=1.8 NRD=16.7056 NRS=1.7533 M=1 R=7.46667
+ SA=75003.1 SB=75003.7 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_89_172#_M1015_g N_Y_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.4424 AS=0.3808 PD=1.91 PS=1.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.9 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g N_VPWR_M1015_d VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.4424 PD=1.42 PS=1.91 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75004.8
+ SB=75001.9 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1007_d N_B_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=1.7472 PD=1.42 PS=5.36 NRD=1.7533 NRS=38.6908 M=1 R=7.46667 SA=75005.3
+ SB=75001.5 A=0.168 P=2.54 MULT=1
DX21_noxref VNB VPB NWDIODE A=14.9916 P=19.84
c_100 VPB 0 1.70138e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__nand3b_4.pxi.spice"
*
.ends
*
*
