* File: sky130_fd_sc_hs__o31ai_4.pxi.spice
* Created: Tue Sep  1 20:18:26 2020
* 
x_PM_SKY130_FD_SC_HS__O31AI_4%A1 N_A1_M1000_g N_A1_c_140_n N_A1_M1011_g
+ N_A1_c_141_n N_A1_M1012_g N_A1_M1004_g N_A1_c_142_n N_A1_M1013_g N_A1_M1022_g
+ N_A1_c_134_n N_A1_c_135_n N_A1_c_136_n N_A1_c_145_n N_A1_M1014_g N_A1_M1029_g
+ N_A1_c_138_n A1 A1 A1 A1 PM_SKY130_FD_SC_HS__O31AI_4%A1
x_PM_SKY130_FD_SC_HS__O31AI_4%A2 N_A2_M1001_g N_A2_c_214_n N_A2_M1010_g
+ N_A2_c_215_n N_A2_c_224_n N_A2_M1015_g N_A2_M1002_g N_A2_c_225_n N_A2_M1016_g
+ N_A2_M1005_g N_A2_c_218_n N_A2_c_219_n N_A2_M1020_g N_A2_c_221_n N_A2_M1017_g
+ A2 A2 A2 PM_SKY130_FD_SC_HS__O31AI_4%A2
x_PM_SKY130_FD_SC_HS__O31AI_4%A3 N_A3_M1006_g N_A3_c_307_n N_A3_c_308_n
+ N_A3_c_316_n N_A3_M1003_g N_A3_M1019_g N_A3_c_317_n N_A3_M1007_g N_A3_M1023_g
+ N_A3_c_318_n N_A3_M1009_g N_A3_c_311_n N_A3_c_312_n N_A3_M1026_g N_A3_c_314_n
+ N_A3_M1027_g A3 A3 A3 PM_SKY130_FD_SC_HS__O31AI_4%A3
x_PM_SKY130_FD_SC_HS__O31AI_4%B1 N_B1_M1018_g N_B1_c_413_n N_B1_M1008_g
+ N_B1_M1021_g N_B1_M1024_g N_B1_c_407_n N_B1_c_408_n N_B1_c_409_n N_B1_c_410_n
+ N_B1_c_416_n N_B1_M1028_g N_B1_c_411_n N_B1_M1025_g B1 B1 B1 N_B1_c_412_n
+ PM_SKY130_FD_SC_HS__O31AI_4%B1
x_PM_SKY130_FD_SC_HS__O31AI_4%A_28_368# N_A_28_368#_M1011_d N_A_28_368#_M1012_d
+ N_A_28_368#_M1014_d N_A_28_368#_M1015_s N_A_28_368#_M1017_s
+ N_A_28_368#_c_472_n N_A_28_368#_c_473_n N_A_28_368#_c_480_n
+ N_A_28_368#_c_474_n N_A_28_368#_c_486_n N_A_28_368#_c_475_n
+ N_A_28_368#_c_498_n N_A_28_368#_c_503_n N_A_28_368#_c_506_n
+ N_A_28_368#_c_507_n N_A_28_368#_c_492_n N_A_28_368#_c_476_n
+ N_A_28_368#_c_514_n N_A_28_368#_c_477_n PM_SKY130_FD_SC_HS__O31AI_4%A_28_368#
x_PM_SKY130_FD_SC_HS__O31AI_4%VPWR N_VPWR_M1011_s N_VPWR_M1013_s N_VPWR_M1008_d
+ N_VPWR_c_550_n N_VPWR_c_551_n VPWR N_VPWR_c_552_n N_VPWR_c_553_n
+ N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_549_n N_VPWR_c_557_n N_VPWR_c_558_n
+ N_VPWR_c_559_n PM_SKY130_FD_SC_HS__O31AI_4%VPWR
x_PM_SKY130_FD_SC_HS__O31AI_4%A_487_368# N_A_487_368#_M1010_d
+ N_A_487_368#_M1016_d N_A_487_368#_M1003_s N_A_487_368#_M1009_s
+ N_A_487_368#_c_639_n N_A_487_368#_c_633_n N_A_487_368#_c_634_n
+ N_A_487_368#_c_635_n N_A_487_368#_c_648_n N_A_487_368#_c_636_n
+ N_A_487_368#_c_652_n N_A_487_368#_c_637_n N_A_487_368#_c_638_n
+ PM_SKY130_FD_SC_HS__O31AI_4%A_487_368#
x_PM_SKY130_FD_SC_HS__O31AI_4%Y N_Y_M1018_d N_Y_M1024_d N_Y_M1003_d N_Y_M1007_d
+ N_Y_M1027_d N_Y_M1028_s N_Y_c_692_n N_Y_c_713_n N_Y_c_697_n N_Y_c_714_n
+ N_Y_c_693_n N_Y_c_723_n N_Y_c_699_n N_Y_c_744_n N_Y_c_694_n N_Y_c_695_n
+ N_Y_c_700_n N_Y_c_701_n N_Y_c_729_n N_Y_c_758_n N_Y_c_696_n Y
+ PM_SKY130_FD_SC_HS__O31AI_4%Y
x_PM_SKY130_FD_SC_HS__O31AI_4%A_27_82# N_A_27_82#_M1000_s N_A_27_82#_M1004_s
+ N_A_27_82#_M1029_s N_A_27_82#_M1002_s N_A_27_82#_M1020_s N_A_27_82#_M1019_d
+ N_A_27_82#_M1026_d N_A_27_82#_M1021_s N_A_27_82#_M1025_s N_A_27_82#_c_808_n
+ N_A_27_82#_c_809_n N_A_27_82#_c_810_n N_A_27_82#_c_811_n N_A_27_82#_c_812_n
+ N_A_27_82#_c_813_n N_A_27_82#_c_814_n N_A_27_82#_c_815_n N_A_27_82#_c_855_n
+ N_A_27_82#_c_816_n N_A_27_82#_c_817_n N_A_27_82#_c_818_n N_A_27_82#_c_819_n
+ N_A_27_82#_c_857_n N_A_27_82#_c_820_n N_A_27_82#_c_821_n N_A_27_82#_c_822_n
+ N_A_27_82#_c_823_n PM_SKY130_FD_SC_HS__O31AI_4%A_27_82#
x_PM_SKY130_FD_SC_HS__O31AI_4%VGND N_VGND_M1000_d N_VGND_M1022_d N_VGND_M1001_d
+ N_VGND_M1005_d N_VGND_M1006_s N_VGND_M1023_s N_VGND_c_938_n N_VGND_c_939_n
+ N_VGND_c_940_n N_VGND_c_941_n N_VGND_c_942_n N_VGND_c_943_n N_VGND_c_944_n
+ VGND N_VGND_c_945_n N_VGND_c_946_n N_VGND_c_947_n N_VGND_c_948_n
+ N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n N_VGND_c_952_n N_VGND_c_953_n
+ N_VGND_c_954_n N_VGND_c_955_n PM_SKY130_FD_SC_HS__O31AI_4%VGND
cc_1 VNB N_A1_M1000_g 0.0301668f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.78
cc_2 VNB N_A1_M1004_g 0.020773f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.78
cc_3 VNB N_A1_M1022_g 0.020773f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.78
cc_4 VNB N_A1_c_134_n 0.0129785f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.425
cc_5 VNB N_A1_c_135_n 0.0532559f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=1.425
cc_6 VNB N_A1_c_136_n 0.00900051f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.675
cc_7 VNB N_A1_M1029_g 0.0216395f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.78
cc_8 VNB N_A1_c_138_n 0.0058476f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.425
cc_9 VNB A1 0.0183603f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_10 VNB N_A2_M1001_g 0.0240055f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.78
cc_11 VNB N_A2_c_214_n 0.0142998f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.765
cc_12 VNB N_A2_c_215_n 0.0125906f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.765
cc_13 VNB N_A2_M1002_g 0.0244227f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.765
cc_14 VNB N_A2_M1005_g 0.0207818f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.425
cc_15 VNB N_A2_c_218_n 0.00622506f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.5
cc_16 VNB N_A2_c_219_n 0.0481464f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.675
cc_17 VNB N_A2_M1020_g 0.0299754f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_18 VNB N_A2_c_221_n 0.00596067f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.78
cc_19 VNB A2 0.00428973f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_20 VNB N_A3_M1006_g 0.0239058f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.78
cc_21 VNB N_A3_c_307_n 0.018252f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.765
cc_22 VNB N_A3_c_308_n 0.00921229f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_23 VNB N_A3_M1019_g 0.0235612f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.78
cc_24 VNB N_A3_M1023_g 0.0222692f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.78
cc_25 VNB N_A3_c_311_n 0.0159079f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.5
cc_26 VNB N_A3_c_312_n 0.0608485f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.675
cc_27 VNB N_A3_M1026_g 0.0295535f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_28 VNB N_A3_c_314_n 0.00622476f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.78
cc_29 VNB A3 0.00465015f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_30 VNB N_B1_M1018_g 0.0207003f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.78
cc_31 VNB N_B1_M1021_g 0.0202302f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_32 VNB N_B1_M1024_g 0.0202302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B1_c_407_n 0.0138734f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_34 VNB N_B1_c_408_n 0.0441119f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_35 VNB N_B1_c_409_n 0.0214806f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.35
cc_36 VNB N_B1_c_410_n 0.0132531f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.78
cc_37 VNB N_B1_c_411_n 0.0192594f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=1.425
cc_38 VNB N_B1_c_412_n 0.00455633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_549_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_692_n 0.00333871f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.78
cc_41 VNB N_Y_c_693_n 0.00711221f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_42 VNB N_Y_c_694_n 9.23665e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_695_n 0.0111386f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_44 VNB N_Y_c_696_n 0.0163097f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.557
cc_45 VNB N_A_27_82#_c_808_n 0.0229545f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.78
cc_46 VNB N_A_27_82#_c_809_n 0.00914199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_82#_c_810_n 0.0140755f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.425
cc_48 VNB N_A_27_82#_c_811_n 0.0025697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_82#_c_812_n 0.00657842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_82#_c_813_n 0.00298673f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.557
cc_51 VNB N_A_27_82#_c_814_n 0.00962965f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_52 VNB N_A_27_82#_c_815_n 0.0019039f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_53 VNB N_A_27_82#_c_816_n 0.0124141f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.565
cc_54 VNB N_A_27_82#_c_817_n 0.0271534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_82#_c_818_n 0.00467923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_27_82#_c_819_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_82#_c_820_n 0.00255379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_27_82#_c_821_n 0.00253903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_82#_c_822_n 0.0025069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_82#_c_823_n 0.00254299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_938_n 0.00782698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_939_n 0.00782698f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.675
cc_63 VNB N_VGND_c_940_n 0.0148817f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.35
cc_64 VNB N_VGND_c_941_n 0.00542539f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.425
cc_65 VNB N_VGND_c_942_n 0.0179129f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_66 VNB N_VGND_c_943_n 0.0193655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_944_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_945_n 0.0193449f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_69 VNB N_VGND_c_946_n 0.016802f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.557
cc_70 VNB N_VGND_c_947_n 0.0195246f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.557
cc_71 VNB N_VGND_c_948_n 0.0611094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_949_n 0.490819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_950_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_951_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_952_n 0.00894416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_953_n 0.0170483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_954_n 0.0237539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_955_n 0.0171644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VPB N_A1_c_140_n 0.0201401f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_80 VPB N_A1_c_141_n 0.0149968f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_81 VPB N_A1_c_142_n 0.0153778f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_82 VPB N_A1_c_135_n 0.0340961f $X=-0.19 $Y=1.66 $X2=1.5 $Y2=1.425
cc_83 VPB N_A1_c_136_n 7.92498e-19 $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.675
cc_84 VPB N_A1_c_145_n 0.0220223f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.765
cc_85 VPB A1 0.018378f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_86 VPB N_A2_c_214_n 0.0227643f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_87 VPB N_A2_c_224_n 0.0166985f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_88 VPB N_A2_c_225_n 0.0162931f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_89 VPB N_A2_c_218_n 0.0096461f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.5
cc_90 VPB N_A2_c_219_n 0.0318151f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.675
cc_91 VPB N_A2_c_221_n 0.0244739f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.78
cc_92 VPB A2 0.012088f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_93 VPB N_A3_c_316_n 0.0173311f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_94 VPB N_A3_c_317_n 0.014664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A3_c_318_n 0.014664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A3_c_312_n 0.0389449f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.675
cc_97 VPB N_A3_c_314_n 0.0213992f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.78
cc_98 VPB A3 0.00971123f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_99 VPB N_B1_c_413_n 0.0186045f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_100 VPB N_B1_c_408_n 0.0325657f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_101 VPB N_B1_c_410_n 0.00116694f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.78
cc_102 VPB N_B1_c_416_n 0.032015f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.78
cc_103 VPB N_B1_c_412_n 0.0120398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_28_368#_c_472_n 0.00739392f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_105 VPB N_A_28_368#_c_473_n 0.0339313f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.35
cc_106 VPB N_A_28_368#_c_474_n 0.00180921f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.5
cc_107 VPB N_A_28_368#_c_475_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.78
cc_108 VPB N_A_28_368#_c_476_n 0.00485881f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.557
cc_109 VPB N_A_28_368#_c_477_n 0.0035924f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_110 VPB N_VPWR_c_550_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.78
cc_111 VPB N_VPWR_c_551_n 0.00582638f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_112 VPB N_VPWR_c_552_n 0.0181665f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.78
cc_113 VPB N_VPWR_c_553_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.675
cc_114 VPB N_VPWR_c_554_n 0.124156f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.78
cc_115 VPB N_VPWR_c_555_n 0.0191816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_549_n 0.0938928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_557_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.557
cc_118 VPB N_VPWR_c_558_n 0.00608948f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.557
cc_119 VPB N_VPWR_c_559_n 0.0354089f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_120 VPB N_A_487_368#_c_633_n 0.00494392f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_121 VPB N_A_487_368#_c_634_n 0.00387025f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.35
cc_122 VPB N_A_487_368#_c_635_n 0.0176561f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.78
cc_123 VPB N_A_487_368#_c_636_n 0.00475813f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.675
cc_124 VPB N_A_487_368#_c_637_n 0.00216079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_487_368#_c_638_n 0.00171072f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_126 VPB N_Y_c_697_n 0.00683455f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.675
cc_127 VPB N_Y_c_693_n 0.0182503f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=2.4
cc_128 VPB N_Y_c_699_n 0.00289633f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_129 VPB N_Y_c_700_n 0.0183125f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_130 VPB N_Y_c_701_n 0.035396f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.557
cc_131 N_A1_M1029_g N_A2_M1001_g 0.0130961f $X=1.925 $Y=0.78 $X2=0 $Y2=0
cc_132 N_A1_c_136_n N_A2_c_214_n 0.0119762f $X=1.91 $Y=1.675 $X2=0 $Y2=0
cc_133 N_A1_c_145_n N_A2_c_214_n 0.0104776f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A1_c_138_n N_A2_c_214_n 0.0130961f $X=1.91 $Y=1.425 $X2=0 $Y2=0
cc_135 A1 N_A2_c_214_n 7.4406e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A1_c_138_n A2 6.94732e-19 $X=1.91 $Y=1.425 $X2=0 $Y2=0
cc_137 A1 N_A_28_368#_c_472_n 0.021684f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A1_c_140_n N_A_28_368#_c_473_n 0.00634858f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A1_c_140_n N_A_28_368#_c_480_n 0.0126853f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A1_c_141_n N_A_28_368#_c_480_n 0.0126853f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_135_n N_A_28_368#_c_480_n 0.00150499f $X=1.5 $Y=1.425 $X2=0 $Y2=0
cc_142 A1 N_A_28_368#_c_480_n 0.0477183f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A1_c_141_n N_A_28_368#_c_474_n 0.00554978f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A1_c_142_n N_A_28_368#_c_474_n 0.00554978f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A1_c_142_n N_A_28_368#_c_486_n 0.0129585f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A1_c_134_n N_A_28_368#_c_486_n 5.38099e-19 $X=1.82 $Y=1.425 $X2=0 $Y2=0
cc_147 N_A1_c_145_n N_A_28_368#_c_486_n 0.0163732f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_148 A1 N_A_28_368#_c_486_n 0.035986f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A1_c_142_n N_A_28_368#_c_475_n 8.85795e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A1_c_145_n N_A_28_368#_c_475_n 0.0107108f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A1_c_135_n N_A_28_368#_c_492_n 0.00104296f $X=1.5 $Y=1.425 $X2=0 $Y2=0
cc_152 A1 N_A_28_368#_c_492_n 0.0150275f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A1_c_142_n N_A_28_368#_c_476_n 6.04745e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A1_c_145_n N_A_28_368#_c_476_n 0.00392567f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A1_c_140_n N_VPWR_c_550_n 0.0141019f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A1_c_141_n N_VPWR_c_550_n 0.0110266f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A1_c_142_n N_VPWR_c_550_n 5.35985e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A1_c_141_n N_VPWR_c_551_n 5.35985e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A1_c_142_n N_VPWR_c_551_n 0.0109623f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A1_c_145_n N_VPWR_c_551_n 0.0056588f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A1_c_140_n N_VPWR_c_552_n 0.00413917f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A1_c_141_n N_VPWR_c_553_n 0.00413917f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A1_c_142_n N_VPWR_c_553_n 0.00413917f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A1_c_145_n N_VPWR_c_554_n 0.00445602f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A1_c_140_n N_VPWR_c_549_n 0.00821237f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A1_c_141_n N_VPWR_c_549_n 0.00817726f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A1_c_142_n N_VPWR_c_549_n 0.00817726f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A1_c_145_n N_VPWR_c_549_n 0.00857462f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A1_M1000_g N_A_27_82#_c_808_n 0.00880243f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_170 N_A1_M1004_g N_A_27_82#_c_808_n 8.60003e-19 $X=0.995 $Y=0.78 $X2=0 $Y2=0
cc_171 N_A1_M1000_g N_A_27_82#_c_809_n 0.0139765f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_172 N_A1_M1004_g N_A_27_82#_c_809_n 0.015662f $X=0.995 $Y=0.78 $X2=0 $Y2=0
cc_173 N_A1_M1022_g N_A_27_82#_c_809_n 0.015662f $X=1.425 $Y=0.78 $X2=0 $Y2=0
cc_174 N_A1_c_134_n N_A_27_82#_c_809_n 0.00350189f $X=1.82 $Y=1.425 $X2=0 $Y2=0
cc_175 N_A1_c_135_n N_A_27_82#_c_809_n 0.00611445f $X=1.5 $Y=1.425 $X2=0 $Y2=0
cc_176 N_A1_M1029_g N_A_27_82#_c_809_n 0.0178224f $X=1.925 $Y=0.78 $X2=0 $Y2=0
cc_177 A1 N_A_27_82#_c_809_n 0.105188f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A1_M1000_g N_A_27_82#_c_810_n 0.00153871f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_179 A1 N_A_27_82#_c_810_n 0.0286342f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A1_M1022_g N_A_27_82#_c_811_n 8.60003e-19 $X=1.425 $Y=0.78 $X2=0 $Y2=0
cc_181 N_A1_M1029_g N_A_27_82#_c_811_n 0.00812924f $X=1.925 $Y=0.78 $X2=0 $Y2=0
cc_182 N_A1_M1029_g N_A_27_82#_c_818_n 0.00161941f $X=1.925 $Y=0.78 $X2=0 $Y2=0
cc_183 N_A1_M1000_g N_VGND_c_938_n 0.00505959f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_184 N_A1_M1004_g N_VGND_c_938_n 0.0106f $X=0.995 $Y=0.78 $X2=0 $Y2=0
cc_185 N_A1_M1022_g N_VGND_c_938_n 0.0013836f $X=1.425 $Y=0.78 $X2=0 $Y2=0
cc_186 N_A1_M1004_g N_VGND_c_939_n 0.0013836f $X=0.995 $Y=0.78 $X2=0 $Y2=0
cc_187 N_A1_M1022_g N_VGND_c_939_n 0.0106f $X=1.425 $Y=0.78 $X2=0 $Y2=0
cc_188 N_A1_M1029_g N_VGND_c_939_n 0.00505959f $X=1.925 $Y=0.78 $X2=0 $Y2=0
cc_189 N_A1_M1000_g N_VGND_c_945_n 0.00523933f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_190 N_A1_M1004_g N_VGND_c_946_n 0.00455951f $X=0.995 $Y=0.78 $X2=0 $Y2=0
cc_191 N_A1_M1022_g N_VGND_c_946_n 0.00455951f $X=1.425 $Y=0.78 $X2=0 $Y2=0
cc_192 N_A1_M1029_g N_VGND_c_947_n 0.00523933f $X=1.925 $Y=0.78 $X2=0 $Y2=0
cc_193 N_A1_M1000_g N_VGND_c_949_n 0.00533081f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_194 N_A1_M1004_g N_VGND_c_949_n 0.00447788f $X=0.995 $Y=0.78 $X2=0 $Y2=0
cc_195 N_A1_M1022_g N_VGND_c_949_n 0.00447788f $X=1.425 $Y=0.78 $X2=0 $Y2=0
cc_196 N_A1_M1029_g N_VGND_c_949_n 0.00533081f $X=1.925 $Y=0.78 $X2=0 $Y2=0
cc_197 N_A2_M1020_g N_A3_M1006_g 0.0238175f $X=4.025 $Y=0.78 $X2=0 $Y2=0
cc_198 N_A2_c_214_n N_A_28_368#_c_475_n 0.0108246f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A2_c_224_n N_A_28_368#_c_475_n 6.21667e-19 $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A2_c_214_n N_A_28_368#_c_498_n 0.0163732f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A2_c_215_n N_A_28_368#_c_498_n 0.00224673f $X=2.66 $Y=1.425 $X2=0 $Y2=0
cc_202 N_A2_c_224_n N_A_28_368#_c_498_n 0.01579f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A2_c_219_n N_A_28_368#_c_498_n 5.23969e-19 $X=3.67 $Y=1.605 $X2=0 $Y2=0
cc_204 A2 N_A_28_368#_c_498_n 0.0311004f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A2_c_225_n N_A_28_368#_c_503_n 0.00254795f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A2_c_219_n N_A_28_368#_c_503_n 0.00195849f $X=3.67 $Y=1.605 $X2=0 $Y2=0
cc_207 A2 N_A_28_368#_c_503_n 0.0281836f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_208 N_A2_c_225_n N_A_28_368#_c_506_n 0.00594002f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A2_c_225_n N_A_28_368#_c_507_n 0.0137847f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A2_c_218_n N_A_28_368#_c_507_n 0.00468491f $X=3.94 $Y=1.605 $X2=0 $Y2=0
cc_211 N_A2_c_219_n N_A_28_368#_c_507_n 7.15844e-19 $X=3.67 $Y=1.605 $X2=0 $Y2=0
cc_212 N_A2_c_221_n N_A_28_368#_c_507_n 0.0124532f $X=4.03 $Y=1.765 $X2=0 $Y2=0
cc_213 A2 N_A_28_368#_c_507_n 0.0109192f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A2_c_214_n N_A_28_368#_c_476_n 0.00386963f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A2_c_224_n N_A_28_368#_c_476_n 6.04745e-19 $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A2_c_225_n N_A_28_368#_c_514_n 0.0048241f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A2_c_214_n N_VPWR_c_554_n 0.00445602f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A2_c_224_n N_VPWR_c_554_n 0.00278257f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A2_c_225_n N_VPWR_c_554_n 0.00279479f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A2_c_221_n N_VPWR_c_554_n 0.00279479f $X=4.03 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A2_c_214_n N_VPWR_c_549_n 0.00858896f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A2_c_224_n N_VPWR_c_549_n 0.0035632f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A2_c_225_n N_VPWR_c_549_n 0.0035495f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A2_c_221_n N_VPWR_c_549_n 0.00357714f $X=4.03 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A2_c_224_n N_A_487_368#_c_639_n 0.0118094f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A2_c_224_n N_A_487_368#_c_633_n 0.011963f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A2_c_225_n N_A_487_368#_c_633_n 0.00936262f $X=3.58 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A2_c_214_n N_A_487_368#_c_634_n 0.00219733f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A2_c_224_n N_A_487_368#_c_634_n 0.00169686f $X=2.86 $Y=1.765 $X2=0
+ $Y2=0
cc_230 N_A2_c_221_n N_A_487_368#_c_635_n 0.0101616f $X=4.03 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A2_c_225_n N_A_487_368#_c_637_n 0.0100612f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A2_c_221_n N_A_487_368#_c_637_n 0.0098754f $X=4.03 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A2_M1020_g N_Y_c_692_n 0.00303574f $X=4.025 $Y=0.78 $X2=0 $Y2=0
cc_234 N_A2_c_221_n N_Y_c_697_n 0.00511995f $X=4.03 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A2_c_225_n N_Y_c_693_n 0.00182693f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A2_c_221_n N_Y_c_693_n 0.0356689f $X=4.03 $Y=1.765 $X2=0 $Y2=0
cc_237 A2 N_Y_c_693_n 0.0146639f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_238 N_A2_M1001_g N_A_27_82#_c_811_n 0.0107656f $X=2.355 $Y=0.78 $X2=0 $Y2=0
cc_239 N_A2_M1001_g N_A_27_82#_c_812_n 0.0162338f $X=2.355 $Y=0.78 $X2=0 $Y2=0
cc_240 N_A2_c_215_n N_A_27_82#_c_812_n 0.00937268f $X=2.66 $Y=1.425 $X2=0 $Y2=0
cc_241 N_A2_M1002_g N_A_27_82#_c_812_n 0.0124466f $X=3.095 $Y=0.78 $X2=0 $Y2=0
cc_242 A2 N_A_27_82#_c_812_n 0.047019f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_243 N_A2_M1002_g N_A_27_82#_c_813_n 0.0146388f $X=3.095 $Y=0.78 $X2=0 $Y2=0
cc_244 N_A2_M1005_g N_A_27_82#_c_813_n 0.00329489f $X=3.595 $Y=0.78 $X2=0 $Y2=0
cc_245 N_A2_M1005_g N_A_27_82#_c_814_n 0.0146865f $X=3.595 $Y=0.78 $X2=0 $Y2=0
cc_246 N_A2_c_218_n N_A_27_82#_c_814_n 0.00282714f $X=3.94 $Y=1.605 $X2=0 $Y2=0
cc_247 N_A2_M1020_g N_A_27_82#_c_814_n 0.0139548f $X=4.025 $Y=0.78 $X2=0 $Y2=0
cc_248 A2 N_A_27_82#_c_814_n 0.0180037f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_249 N_A2_M1001_g N_A_27_82#_c_818_n 0.00580256f $X=2.355 $Y=0.78 $X2=0 $Y2=0
cc_250 N_A2_c_214_n N_A_27_82#_c_818_n 2.37425e-19 $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A2_M1002_g N_A_27_82#_c_819_n 0.00116367f $X=3.095 $Y=0.78 $X2=0 $Y2=0
cc_252 N_A2_c_219_n N_A_27_82#_c_819_n 0.00396026f $X=3.67 $Y=1.605 $X2=0 $Y2=0
cc_253 A2 N_A_27_82#_c_819_n 0.0282341f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_254 N_A2_M1001_g N_VGND_c_940_n 0.00828548f $X=2.355 $Y=0.78 $X2=0 $Y2=0
cc_255 N_A2_M1002_g N_VGND_c_940_n 0.00831784f $X=3.095 $Y=0.78 $X2=0 $Y2=0
cc_256 N_A2_M1002_g N_VGND_c_941_n 6.63069e-19 $X=3.095 $Y=0.78 $X2=0 $Y2=0
cc_257 N_A2_M1005_g N_VGND_c_941_n 0.00972691f $X=3.595 $Y=0.78 $X2=0 $Y2=0
cc_258 N_A2_M1020_g N_VGND_c_941_n 0.00969098f $X=4.025 $Y=0.78 $X2=0 $Y2=0
cc_259 N_A2_M1002_g N_VGND_c_943_n 0.00523933f $X=3.095 $Y=0.78 $X2=0 $Y2=0
cc_260 N_A2_M1005_g N_VGND_c_943_n 0.00455951f $X=3.595 $Y=0.78 $X2=0 $Y2=0
cc_261 N_A2_M1001_g N_VGND_c_947_n 0.00523933f $X=2.355 $Y=0.78 $X2=0 $Y2=0
cc_262 N_A2_M1001_g N_VGND_c_949_n 0.00533081f $X=2.355 $Y=0.78 $X2=0 $Y2=0
cc_263 N_A2_M1002_g N_VGND_c_949_n 0.00533081f $X=3.095 $Y=0.78 $X2=0 $Y2=0
cc_264 N_A2_M1005_g N_VGND_c_949_n 0.00447788f $X=3.595 $Y=0.78 $X2=0 $Y2=0
cc_265 N_A2_M1020_g N_VGND_c_949_n 0.00447788f $X=4.025 $Y=0.78 $X2=0 $Y2=0
cc_266 N_A2_M1020_g N_VGND_c_953_n 0.00455951f $X=4.025 $Y=0.78 $X2=0 $Y2=0
cc_267 N_A3_M1026_g N_B1_M1018_g 0.0235058f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_268 N_A3_c_314_n N_B1_c_413_n 0.0244665f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_269 N_A3_c_314_n N_B1_c_408_n 0.0289705f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_270 N_A3_c_312_n N_B1_c_412_n 2.75683e-19 $X=6.08 $Y=1.555 $X2=0 $Y2=0
cc_271 N_A3_M1026_g N_B1_c_412_n 0.00590426f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_272 N_A3_c_314_n N_B1_c_412_n 0.0136806f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_273 A3 N_B1_c_412_n 0.0277795f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_274 N_A3_c_316_n N_VPWR_c_554_n 0.00278257f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_275 N_A3_c_317_n N_VPWR_c_554_n 0.00278271f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_276 N_A3_c_318_n N_VPWR_c_554_n 0.00278271f $X=5.99 $Y=1.765 $X2=0 $Y2=0
cc_277 N_A3_c_314_n N_VPWR_c_554_n 0.0044313f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_278 N_A3_c_316_n N_VPWR_c_549_n 0.00358623f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_279 N_A3_c_317_n N_VPWR_c_549_n 0.00353823f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A3_c_318_n N_VPWR_c_549_n 0.00353823f $X=5.99 $Y=1.765 $X2=0 $Y2=0
cc_281 N_A3_c_314_n N_VPWR_c_549_n 0.00854637f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_282 N_A3_c_316_n N_A_487_368#_c_635_n 0.012762f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_283 N_A3_c_316_n N_A_487_368#_c_648_n 0.0117018f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_284 N_A3_c_317_n N_A_487_368#_c_636_n 0.0128349f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A3_c_318_n N_A_487_368#_c_636_n 0.0128349f $X=5.99 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A3_c_314_n N_A_487_368#_c_636_n 0.00408436f $X=6.44 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_A3_c_314_n N_A_487_368#_c_652_n 0.00604065f $X=6.44 $Y=1.765 $X2=0
+ $Y2=0
cc_288 N_A3_c_316_n N_A_487_368#_c_638_n 0.00175197f $X=5.09 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_A3_M1006_g N_Y_c_692_n 0.0058695f $X=4.455 $Y=0.78 $X2=0 $Y2=0
cc_290 N_A3_c_307_n N_Y_c_692_n 0.00795652f $X=4.835 $Y=1.425 $X2=0 $Y2=0
cc_291 N_A3_c_308_n N_Y_c_692_n 0.00348927f $X=4.53 $Y=1.425 $X2=0 $Y2=0
cc_292 N_A3_M1019_g N_Y_c_692_n 0.00350741f $X=5.395 $Y=0.78 $X2=0 $Y2=0
cc_293 N_A3_c_312_n N_Y_c_692_n 3.45584e-19 $X=6.08 $Y=1.555 $X2=0 $Y2=0
cc_294 A3 N_Y_c_692_n 0.0153081f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_295 N_A3_M1006_g N_Y_c_713_n 0.00644113f $X=4.455 $Y=0.78 $X2=0 $Y2=0
cc_296 N_A3_c_316_n N_Y_c_714_n 0.0126853f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_297 N_A3_c_317_n N_Y_c_714_n 0.0120074f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_298 N_A3_c_312_n N_Y_c_714_n 0.00130507f $X=6.08 $Y=1.555 $X2=0 $Y2=0
cc_299 A3 N_Y_c_714_n 0.042432f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_300 N_A3_c_307_n N_Y_c_693_n 0.00503033f $X=4.835 $Y=1.425 $X2=0 $Y2=0
cc_301 N_A3_c_308_n N_Y_c_693_n 0.00621365f $X=4.53 $Y=1.425 $X2=0 $Y2=0
cc_302 N_A3_c_316_n N_Y_c_693_n 0.0043164f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_303 N_A3_c_312_n N_Y_c_693_n 0.00227395f $X=6.08 $Y=1.555 $X2=0 $Y2=0
cc_304 A3 N_Y_c_693_n 0.0323075f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_305 N_A3_c_318_n N_Y_c_723_n 0.0120074f $X=5.99 $Y=1.765 $X2=0 $Y2=0
cc_306 N_A3_c_311_n N_Y_c_723_n 0.0066691f $X=6.35 $Y=1.555 $X2=0 $Y2=0
cc_307 N_A3_c_314_n N_Y_c_723_n 0.0150982f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_308 A3 N_Y_c_723_n 0.0119829f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_309 N_A3_c_314_n N_Y_c_699_n 0.00464012f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_310 N_A3_M1026_g N_Y_c_694_n 4.30079e-19 $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_311 N_A3_c_316_n N_Y_c_729_n 4.46973e-19 $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_312 N_A3_c_317_n N_Y_c_729_n 0.00907138f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A3_c_318_n N_Y_c_729_n 0.00904709f $X=5.99 $Y=1.765 $X2=0 $Y2=0
cc_314 N_A3_c_312_n N_Y_c_729_n 0.00143667f $X=6.08 $Y=1.555 $X2=0 $Y2=0
cc_315 N_A3_c_314_n N_Y_c_729_n 4.45174e-19 $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_316 A3 N_Y_c_729_n 0.0237598f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_317 N_A3_c_307_n N_Y_c_696_n 0.0152657f $X=4.835 $Y=1.425 $X2=0 $Y2=0
cc_318 N_A3_M1019_g N_Y_c_696_n 0.0125331f $X=5.395 $Y=0.78 $X2=0 $Y2=0
cc_319 N_A3_M1023_g N_Y_c_696_n 0.011771f $X=5.825 $Y=0.78 $X2=0 $Y2=0
cc_320 N_A3_c_311_n N_Y_c_696_n 0.00432054f $X=6.35 $Y=1.555 $X2=0 $Y2=0
cc_321 N_A3_c_312_n N_Y_c_696_n 0.00310668f $X=6.08 $Y=1.555 $X2=0 $Y2=0
cc_322 N_A3_M1026_g N_Y_c_696_n 0.012224f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_323 A3 N_Y_c_696_n 0.0979855f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_324 N_A3_M1006_g N_A_27_82#_c_814_n 2.37852e-19 $X=4.455 $Y=0.78 $X2=0 $Y2=0
cc_325 N_A3_M1023_g N_A_27_82#_c_855_n 0.00930211f $X=5.825 $Y=0.78 $X2=0 $Y2=0
cc_326 N_A3_M1026_g N_A_27_82#_c_855_n 0.00985212f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_327 N_A3_M1006_g N_A_27_82#_c_857_n 0.0156099f $X=4.455 $Y=0.78 $X2=0 $Y2=0
cc_328 N_A3_c_307_n N_A_27_82#_c_857_n 8.27297e-19 $X=4.835 $Y=1.425 $X2=0 $Y2=0
cc_329 N_A3_M1019_g N_A_27_82#_c_857_n 0.0104597f $X=5.395 $Y=0.78 $X2=0 $Y2=0
cc_330 N_A3_M1019_g N_A_27_82#_c_820_n 0.0106333f $X=5.395 $Y=0.78 $X2=0 $Y2=0
cc_331 N_A3_M1023_g N_A_27_82#_c_820_n 0.00747156f $X=5.825 $Y=0.78 $X2=0 $Y2=0
cc_332 N_A3_M1026_g N_A_27_82#_c_820_n 0.00116516f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_333 N_A3_M1023_g N_A_27_82#_c_821_n 8.49064e-19 $X=5.825 $Y=0.78 $X2=0 $Y2=0
cc_334 N_A3_M1026_g N_A_27_82#_c_821_n 0.00553413f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_335 N_A3_M1006_g N_VGND_c_941_n 4.95268e-19 $X=4.455 $Y=0.78 $X2=0 $Y2=0
cc_336 N_A3_M1019_g N_VGND_c_942_n 0.00418922f $X=5.395 $Y=0.78 $X2=0 $Y2=0
cc_337 N_A3_M1023_g N_VGND_c_942_n 0.00411482f $X=5.825 $Y=0.78 $X2=0 $Y2=0
cc_338 N_A3_M1026_g N_VGND_c_948_n 0.00412495f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_339 N_A3_M1006_g N_VGND_c_949_n 0.00533081f $X=4.455 $Y=0.78 $X2=0 $Y2=0
cc_340 N_A3_M1019_g N_VGND_c_949_n 0.00533081f $X=5.395 $Y=0.78 $X2=0 $Y2=0
cc_341 N_A3_M1023_g N_VGND_c_949_n 0.00533081f $X=5.825 $Y=0.78 $X2=0 $Y2=0
cc_342 N_A3_M1026_g N_VGND_c_949_n 0.00533081f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_343 N_A3_M1006_g N_VGND_c_953_n 0.0042391f $X=4.455 $Y=0.78 $X2=0 $Y2=0
cc_344 N_A3_M1006_g N_VGND_c_954_n 0.00555179f $X=4.455 $Y=0.78 $X2=0 $Y2=0
cc_345 N_A3_M1019_g N_VGND_c_954_n 0.00727635f $X=5.395 $Y=0.78 $X2=0 $Y2=0
cc_346 N_A3_M1023_g N_VGND_c_955_n 0.00344286f $X=5.825 $Y=0.78 $X2=0 $Y2=0
cc_347 N_A3_M1026_g N_VGND_c_955_n 0.00342357f $X=6.425 $Y=0.78 $X2=0 $Y2=0
cc_348 N_B1_c_413_n N_VPWR_c_554_n 0.00445602f $X=6.94 $Y=1.765 $X2=0 $Y2=0
cc_349 N_B1_c_416_n N_VPWR_c_555_n 0.00445602f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_350 N_B1_c_413_n N_VPWR_c_549_n 0.00862233f $X=6.94 $Y=1.765 $X2=0 $Y2=0
cc_351 N_B1_c_416_n N_VPWR_c_549_n 0.00865213f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_352 N_B1_c_413_n N_VPWR_c_559_n 0.00420542f $X=6.94 $Y=1.765 $X2=0 $Y2=0
cc_353 N_B1_c_416_n N_VPWR_c_559_n 0.00565407f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_354 N_B1_c_413_n N_A_487_368#_c_636_n 3.17734e-19 $X=6.94 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_B1_c_412_n N_Y_c_723_n 0.0124612f $X=7.625 $Y=1.515 $X2=0 $Y2=0
cc_356 N_B1_c_413_n N_Y_c_699_n 0.0144328f $X=6.94 $Y=1.765 $X2=0 $Y2=0
cc_357 N_B1_c_413_n N_Y_c_744_n 0.0139279f $X=6.94 $Y=1.765 $X2=0 $Y2=0
cc_358 N_B1_c_407_n N_Y_c_744_n 0.00676058f $X=8.045 $Y=1.425 $X2=0 $Y2=0
cc_359 N_B1_c_408_n N_Y_c_744_n 0.00402819f $X=7.79 $Y=1.425 $X2=0 $Y2=0
cc_360 N_B1_c_416_n N_Y_c_744_n 0.0180205f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_361 N_B1_c_412_n N_Y_c_744_n 0.0694754f $X=7.625 $Y=1.515 $X2=0 $Y2=0
cc_362 N_B1_M1018_g N_Y_c_694_n 0.003332f $X=6.855 $Y=0.78 $X2=0 $Y2=0
cc_363 N_B1_c_408_n N_Y_c_694_n 0.00227305f $X=7.79 $Y=1.425 $X2=0 $Y2=0
cc_364 N_B1_M1021_g N_Y_c_695_n 0.012086f $X=7.285 $Y=0.78 $X2=0 $Y2=0
cc_365 N_B1_M1024_g N_Y_c_695_n 0.012086f $X=7.715 $Y=0.78 $X2=0 $Y2=0
cc_366 N_B1_c_407_n N_Y_c_695_n 0.00360194f $X=8.045 $Y=1.425 $X2=0 $Y2=0
cc_367 N_B1_c_408_n N_Y_c_695_n 0.00226461f $X=7.79 $Y=1.425 $X2=0 $Y2=0
cc_368 N_B1_c_411_n N_Y_c_695_n 0.0050901f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_369 N_B1_c_416_n N_Y_c_700_n 0.00774852f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_370 N_B1_c_416_n N_Y_c_701_n 0.0156099f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_371 N_B1_c_413_n N_Y_c_758_n 4.27055e-19 $X=6.94 $Y=1.765 $X2=0 $Y2=0
cc_372 N_B1_c_408_n N_Y_c_758_n 3.21196e-19 $X=7.79 $Y=1.425 $X2=0 $Y2=0
cc_373 N_B1_c_412_n N_Y_c_758_n 0.0254782f $X=7.625 $Y=1.515 $X2=0 $Y2=0
cc_374 N_B1_M1018_g N_Y_c_696_n 0.00834439f $X=6.855 $Y=0.78 $X2=0 $Y2=0
cc_375 N_B1_c_412_n N_Y_c_696_n 0.110395f $X=7.625 $Y=1.515 $X2=0 $Y2=0
cc_376 N_B1_M1024_g N_A_27_82#_c_816_n 0.00787355f $X=7.715 $Y=0.78 $X2=0 $Y2=0
cc_377 N_B1_c_411_n N_A_27_82#_c_816_n 0.0123592f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_378 N_B1_c_411_n N_A_27_82#_c_817_n 0.00131802f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_379 N_B1_M1018_g N_A_27_82#_c_821_n 0.00506303f $X=6.855 $Y=0.78 $X2=0 $Y2=0
cc_380 N_B1_M1021_g N_A_27_82#_c_821_n 6.42481e-19 $X=7.285 $Y=0.78 $X2=0 $Y2=0
cc_381 N_B1_M1018_g N_A_27_82#_c_822_n 0.00869307f $X=6.855 $Y=0.78 $X2=0 $Y2=0
cc_382 N_B1_M1021_g N_A_27_82#_c_822_n 0.00787355f $X=7.285 $Y=0.78 $X2=0 $Y2=0
cc_383 N_B1_M1018_g N_A_27_82#_c_823_n 5.57235e-19 $X=6.855 $Y=0.78 $X2=0 $Y2=0
cc_384 N_B1_M1021_g N_A_27_82#_c_823_n 0.00451712f $X=7.285 $Y=0.78 $X2=0 $Y2=0
cc_385 N_B1_M1024_g N_A_27_82#_c_823_n 0.00472539f $X=7.715 $Y=0.78 $X2=0 $Y2=0
cc_386 N_B1_c_411_n N_A_27_82#_c_823_n 5.73274e-19 $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_387 N_B1_M1018_g N_VGND_c_948_n 0.00394994f $X=6.855 $Y=0.78 $X2=0 $Y2=0
cc_388 N_B1_M1021_g N_VGND_c_948_n 0.00393982f $X=7.285 $Y=0.78 $X2=0 $Y2=0
cc_389 N_B1_M1024_g N_VGND_c_948_n 0.00393982f $X=7.715 $Y=0.78 $X2=0 $Y2=0
cc_390 N_B1_c_411_n N_VGND_c_948_n 0.00393982f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_391 N_B1_M1018_g N_VGND_c_949_n 0.00533081f $X=6.855 $Y=0.78 $X2=0 $Y2=0
cc_392 N_B1_M1021_g N_VGND_c_949_n 0.00533081f $X=7.285 $Y=0.78 $X2=0 $Y2=0
cc_393 N_B1_M1024_g N_VGND_c_949_n 0.00533081f $X=7.715 $Y=0.78 $X2=0 $Y2=0
cc_394 N_B1_c_411_n N_VGND_c_949_n 0.00533081f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_395 N_A_28_368#_c_480_n N_VPWR_M1011_s 0.00359365f $X=1.1 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_396 N_A_28_368#_c_486_n N_VPWR_M1013_s 0.00483578f $X=1.97 $Y=2.035 $X2=0
+ $Y2=0
cc_397 N_A_28_368#_c_473_n N_VPWR_c_550_n 0.0462948f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_398 N_A_28_368#_c_480_n N_VPWR_c_550_n 0.0171813f $X=1.1 $Y=2.035 $X2=0 $Y2=0
cc_399 N_A_28_368#_c_474_n N_VPWR_c_550_n 0.0449718f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_400 N_A_28_368#_c_474_n N_VPWR_c_551_n 0.0449718f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_401 N_A_28_368#_c_486_n N_VPWR_c_551_n 0.0202249f $X=1.97 $Y=2.035 $X2=0
+ $Y2=0
cc_402 N_A_28_368#_c_475_n N_VPWR_c_551_n 0.0266809f $X=2.135 $Y=2.815 $X2=0
+ $Y2=0
cc_403 N_A_28_368#_c_473_n N_VPWR_c_552_n 0.011066f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_404 N_A_28_368#_c_474_n N_VPWR_c_553_n 0.00749631f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_405 N_A_28_368#_c_475_n N_VPWR_c_554_n 0.014552f $X=2.135 $Y=2.815 $X2=0
+ $Y2=0
cc_406 N_A_28_368#_c_473_n N_VPWR_c_549_n 0.00915947f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_407 N_A_28_368#_c_474_n N_VPWR_c_549_n 0.0062048f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_408 N_A_28_368#_c_475_n N_VPWR_c_549_n 0.0119791f $X=2.135 $Y=2.815 $X2=0
+ $Y2=0
cc_409 N_A_28_368#_c_507_n N_VPWR_c_549_n 0.00194189f $X=4.14 $Y=2.455 $X2=0
+ $Y2=0
cc_410 N_A_28_368#_c_498_n N_A_487_368#_M1010_d 0.00484339f $X=2.97 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_411 N_A_28_368#_c_507_n N_A_487_368#_M1016_d 0.00523323f $X=4.14 $Y=2.455
+ $X2=0 $Y2=0
cc_412 N_A_28_368#_c_498_n N_A_487_368#_c_639_n 0.0202249f $X=2.97 $Y=2.035
+ $X2=0 $Y2=0
cc_413 N_A_28_368#_M1015_s N_A_487_368#_c_633_n 0.00615455f $X=2.935 $Y=1.84
+ $X2=0 $Y2=0
cc_414 N_A_28_368#_c_507_n N_A_487_368#_c_633_n 0.0096007f $X=4.14 $Y=2.455
+ $X2=0 $Y2=0
cc_415 N_A_28_368#_c_514_n N_A_487_368#_c_633_n 0.0233667f $X=3.135 $Y=2.455
+ $X2=0 $Y2=0
cc_416 N_A_28_368#_c_475_n N_A_487_368#_c_634_n 0.00371331f $X=2.135 $Y=2.815
+ $X2=0 $Y2=0
cc_417 N_A_28_368#_M1017_s N_A_487_368#_c_635_n 0.00355467f $X=4.105 $Y=1.84
+ $X2=0 $Y2=0
cc_418 N_A_28_368#_c_507_n N_A_487_368#_c_635_n 0.00429117f $X=4.14 $Y=2.455
+ $X2=0 $Y2=0
cc_419 N_A_28_368#_c_477_n N_A_487_368#_c_635_n 0.0223455f $X=4.305 $Y=2.455
+ $X2=0 $Y2=0
cc_420 N_A_28_368#_c_507_n N_A_487_368#_c_637_n 0.0158897f $X=4.14 $Y=2.455
+ $X2=0 $Y2=0
cc_421 N_A_28_368#_c_514_n N_A_487_368#_c_637_n 0.00114028f $X=3.135 $Y=2.455
+ $X2=0 $Y2=0
cc_422 N_A_28_368#_c_477_n N_Y_c_697_n 0.0242398f $X=4.305 $Y=2.455 $X2=0 $Y2=0
cc_423 N_A_28_368#_M1017_s N_Y_c_693_n 0.00638842f $X=4.105 $Y=1.84 $X2=0 $Y2=0
cc_424 N_A_28_368#_c_503_n N_Y_c_693_n 0.00498715f $X=3.135 $Y=2.12 $X2=0 $Y2=0
cc_425 N_A_28_368#_c_506_n N_Y_c_693_n 8.15755e-19 $X=3.135 $Y=2.37 $X2=0 $Y2=0
cc_426 N_A_28_368#_c_507_n N_Y_c_693_n 0.00857797f $X=4.14 $Y=2.455 $X2=0 $Y2=0
cc_427 N_A_28_368#_c_477_n N_Y_c_693_n 0.0216785f $X=4.305 $Y=2.455 $X2=0 $Y2=0
cc_428 N_A_28_368#_c_476_n N_A_27_82#_c_818_n 0.0116847f $X=2.135 $Y=1.985 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_554_n N_A_487_368#_c_633_n 0.0532992f $X=7.05 $Y=3.33 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_549_n N_A_487_368#_c_633_n 0.0303501f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_431 N_VPWR_c_551_n N_A_487_368#_c_634_n 0.00314404f $X=1.635 $Y=2.455 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_554_n N_A_487_368#_c_634_n 0.0236039f $X=7.05 $Y=3.33 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_549_n N_A_487_368#_c_634_n 0.012761f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_554_n N_A_487_368#_c_635_n 0.0752014f $X=7.05 $Y=3.33 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_549_n N_A_487_368#_c_635_n 0.0431333f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_436 N_VPWR_c_554_n N_A_487_368#_c_636_n 0.0639627f $X=7.05 $Y=3.33 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_549_n N_A_487_368#_c_636_n 0.035724f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_438 N_VPWR_c_559_n N_A_487_368#_c_636_n 0.00292455f $X=7.165 $Y=2.455 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_554_n N_A_487_368#_c_637_n 0.0223621f $X=7.05 $Y=3.33 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_549_n N_A_487_368#_c_637_n 0.0124265f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_441 N_VPWR_c_554_n N_A_487_368#_c_638_n 0.017869f $X=7.05 $Y=3.33 $X2=0 $Y2=0
cc_442 N_VPWR_c_549_n N_A_487_368#_c_638_n 0.00965079f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_554_n N_Y_c_699_n 0.0145938f $X=7.05 $Y=3.33 $X2=0 $Y2=0
cc_444 N_VPWR_c_549_n N_Y_c_699_n 0.0120466f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_445 N_VPWR_c_559_n N_Y_c_699_n 0.0267725f $X=7.165 $Y=2.455 $X2=0 $Y2=0
cc_446 N_VPWR_M1008_d N_Y_c_744_n 0.0256445f $X=7.015 $Y=1.84 $X2=0 $Y2=0
cc_447 N_VPWR_c_559_n N_Y_c_744_n 0.0757448f $X=7.165 $Y=2.455 $X2=0 $Y2=0
cc_448 N_VPWR_c_555_n N_Y_c_701_n 0.0145938f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_449 N_VPWR_c_549_n N_Y_c_701_n 0.0120466f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_450 N_VPWR_c_559_n N_Y_c_701_n 0.0267725f $X=7.165 $Y=2.455 $X2=0 $Y2=0
cc_451 N_A_487_368#_c_635_n N_Y_M1003_d 0.00287371f $X=5.15 $Y=2.99 $X2=0 $Y2=0
cc_452 N_A_487_368#_c_636_n N_Y_M1007_d 0.00197722f $X=6.13 $Y=2.99 $X2=0 $Y2=0
cc_453 N_A_487_368#_c_635_n N_Y_c_697_n 0.019616f $X=5.15 $Y=2.99 $X2=0 $Y2=0
cc_454 N_A_487_368#_M1003_s N_Y_c_714_n 0.00384138f $X=5.165 $Y=1.84 $X2=0 $Y2=0
cc_455 N_A_487_368#_c_648_n N_Y_c_714_n 0.0154248f $X=5.315 $Y=2.455 $X2=0 $Y2=0
cc_456 N_A_487_368#_M1009_s N_Y_c_723_n 0.00465988f $X=6.065 $Y=1.84 $X2=0 $Y2=0
cc_457 N_A_487_368#_c_652_n N_Y_c_723_n 0.0154248f $X=6.215 $Y=2.455 $X2=0 $Y2=0
cc_458 N_A_487_368#_c_636_n N_Y_c_699_n 0.00395311f $X=6.13 $Y=2.99 $X2=0 $Y2=0
cc_459 N_A_487_368#_c_648_n N_Y_c_729_n 0.0298377f $X=5.315 $Y=2.455 $X2=0 $Y2=0
cc_460 N_A_487_368#_c_636_n N_Y_c_729_n 0.0160777f $X=6.13 $Y=2.99 $X2=0 $Y2=0
cc_461 N_A_487_368#_c_652_n N_Y_c_729_n 0.0298377f $X=6.215 $Y=2.455 $X2=0 $Y2=0
cc_462 N_Y_c_696_n N_A_27_82#_M1019_d 0.00176891f $X=6.905 $Y=1.05 $X2=0 $Y2=0
cc_463 N_Y_c_696_n N_A_27_82#_M1026_d 0.00213686f $X=6.905 $Y=1.05 $X2=0 $Y2=0
cc_464 N_Y_c_695_n N_A_27_82#_M1021_s 0.00179223f $X=7.93 $Y=1.005 $X2=0 $Y2=0
cc_465 N_Y_c_713_n N_A_27_82#_c_814_n 0.00855301f $X=4.665 $Y=1.095 $X2=0 $Y2=0
cc_466 N_Y_c_693_n N_A_27_82#_c_814_n 0.0172686f $X=4.97 $Y=2.035 $X2=0 $Y2=0
cc_467 N_Y_c_696_n N_A_27_82#_c_855_n 0.0298909f $X=6.905 $Y=1.05 $X2=0 $Y2=0
cc_468 N_Y_M1024_d N_A_27_82#_c_816_n 0.00252058f $X=7.79 $Y=0.41 $X2=0 $Y2=0
cc_469 N_Y_c_695_n N_A_27_82#_c_816_n 0.0128702f $X=7.93 $Y=1.005 $X2=0 $Y2=0
cc_470 N_Y_c_695_n N_A_27_82#_c_817_n 0.0112546f $X=7.93 $Y=1.005 $X2=0 $Y2=0
cc_471 N_Y_c_700_n N_A_27_82#_c_817_n 0.0094281f $X=8.36 $Y=2.12 $X2=0 $Y2=0
cc_472 N_Y_c_713_n N_A_27_82#_c_857_n 0.0090121f $X=4.665 $Y=1.095 $X2=0 $Y2=0
cc_473 N_Y_c_696_n N_A_27_82#_c_857_n 0.0684999f $X=6.905 $Y=1.05 $X2=0 $Y2=0
cc_474 N_Y_c_696_n N_A_27_82#_c_821_n 0.0117841f $X=6.905 $Y=1.05 $X2=0 $Y2=0
cc_475 N_Y_M1018_d N_A_27_82#_c_822_n 0.00252058f $X=6.93 $Y=0.41 $X2=0 $Y2=0
cc_476 N_Y_c_694_n N_A_27_82#_c_822_n 0.0128479f $X=7.035 $Y=1.05 $X2=0 $Y2=0
cc_477 N_Y_c_696_n N_A_27_82#_c_822_n 0.00306481f $X=6.905 $Y=1.05 $X2=0 $Y2=0
cc_478 N_Y_c_695_n N_A_27_82#_c_823_n 0.0168031f $X=7.93 $Y=1.005 $X2=0 $Y2=0
cc_479 N_Y_c_713_n N_VGND_M1006_s 8.65291e-19 $X=4.665 $Y=1.095 $X2=0 $Y2=0
cc_480 N_Y_c_696_n N_VGND_M1006_s 0.00966998f $X=6.905 $Y=1.05 $X2=0 $Y2=0
cc_481 N_Y_c_696_n N_VGND_M1023_s 0.00502568f $X=6.905 $Y=1.05 $X2=0 $Y2=0
cc_482 N_A_27_82#_c_809_n N_VGND_M1000_d 0.00254178f $X=1.975 $Y=1.05 $X2=-0.19
+ $Y2=-0.245
cc_483 N_A_27_82#_c_809_n N_VGND_M1022_d 0.00254178f $X=1.975 $Y=1.05 $X2=0
+ $Y2=0
cc_484 N_A_27_82#_c_812_n N_VGND_M1001_d 0.00744839f $X=3.145 $Y=1.095 $X2=0
+ $Y2=0
cc_485 N_A_27_82#_c_814_n N_VGND_M1005_d 0.00176461f $X=4.155 $Y=1.095 $X2=0
+ $Y2=0
cc_486 N_A_27_82#_c_857_n N_VGND_M1006_s 0.017452f $X=5.445 $Y=0.615 $X2=0 $Y2=0
cc_487 N_A_27_82#_c_855_n N_VGND_M1023_s 0.00856341f $X=6.475 $Y=0.665 $X2=0
+ $Y2=0
cc_488 N_A_27_82#_c_808_n N_VGND_c_938_n 0.0142986f $X=0.28 $Y=0.555 $X2=0 $Y2=0
cc_489 N_A_27_82#_c_809_n N_VGND_c_938_n 0.0216074f $X=1.975 $Y=1.05 $X2=0 $Y2=0
cc_490 N_A_27_82#_c_809_n N_VGND_c_939_n 0.0216074f $X=1.975 $Y=1.05 $X2=0 $Y2=0
cc_491 N_A_27_82#_c_811_n N_VGND_c_939_n 0.0142986f $X=2.14 $Y=0.555 $X2=0 $Y2=0
cc_492 N_A_27_82#_c_811_n N_VGND_c_940_n 0.0304043f $X=2.14 $Y=0.555 $X2=0 $Y2=0
cc_493 N_A_27_82#_c_812_n N_VGND_c_940_n 0.0327668f $X=3.145 $Y=1.095 $X2=0
+ $Y2=0
cc_494 N_A_27_82#_c_813_n N_VGND_c_940_n 0.0310329f $X=3.31 $Y=0.555 $X2=0 $Y2=0
cc_495 N_A_27_82#_c_813_n N_VGND_c_941_n 0.0176756f $X=3.31 $Y=0.555 $X2=0 $Y2=0
cc_496 N_A_27_82#_c_814_n N_VGND_c_941_n 0.0170777f $X=4.155 $Y=1.095 $X2=0
+ $Y2=0
cc_497 N_A_27_82#_c_815_n N_VGND_c_941_n 0.0107221f $X=4.24 $Y=0.555 $X2=0 $Y2=0
cc_498 N_A_27_82#_c_855_n N_VGND_c_942_n 0.00294479f $X=6.475 $Y=0.665 $X2=0
+ $Y2=0
cc_499 N_A_27_82#_c_857_n N_VGND_c_942_n 0.00236055f $X=5.445 $Y=0.615 $X2=0
+ $Y2=0
cc_500 N_A_27_82#_c_820_n N_VGND_c_942_n 0.0121348f $X=5.775 $Y=0.615 $X2=0
+ $Y2=0
cc_501 N_A_27_82#_c_813_n N_VGND_c_943_n 0.0125377f $X=3.31 $Y=0.555 $X2=0 $Y2=0
cc_502 N_A_27_82#_c_808_n N_VGND_c_945_n 0.0125377f $X=0.28 $Y=0.555 $X2=0 $Y2=0
cc_503 N_A_27_82#_c_811_n N_VGND_c_947_n 0.0124701f $X=2.14 $Y=0.555 $X2=0 $Y2=0
cc_504 N_A_27_82#_c_855_n N_VGND_c_948_n 0.0029521f $X=6.475 $Y=0.665 $X2=0
+ $Y2=0
cc_505 N_A_27_82#_c_816_n N_VGND_c_948_n 0.00999194f $X=8.265 $Y=0.475 $X2=0
+ $Y2=0
cc_506 N_A_27_82#_c_821_n N_VGND_c_948_n 0.0119271f $X=6.64 $Y=0.475 $X2=0 $Y2=0
cc_507 N_A_27_82#_c_822_n N_VGND_c_948_n 0.0500146f $X=7.335 $Y=0.57 $X2=0 $Y2=0
cc_508 N_A_27_82#_c_808_n N_VGND_c_949_n 0.0117961f $X=0.28 $Y=0.555 $X2=0 $Y2=0
cc_509 N_A_27_82#_c_811_n N_VGND_c_949_n 0.0117748f $X=2.14 $Y=0.555 $X2=0 $Y2=0
cc_510 N_A_27_82#_c_813_n N_VGND_c_949_n 0.0117961f $X=3.31 $Y=0.555 $X2=0 $Y2=0
cc_511 N_A_27_82#_c_815_n N_VGND_c_949_n 0.00605288f $X=4.24 $Y=0.555 $X2=0
+ $Y2=0
cc_512 N_A_27_82#_c_855_n N_VGND_c_949_n 0.0122394f $X=6.475 $Y=0.665 $X2=0
+ $Y2=0
cc_513 N_A_27_82#_c_816_n N_VGND_c_949_n 0.00936755f $X=8.265 $Y=0.475 $X2=0
+ $Y2=0
cc_514 N_A_27_82#_c_857_n N_VGND_c_949_n 0.0147815f $X=5.445 $Y=0.615 $X2=0
+ $Y2=0
cc_515 N_A_27_82#_c_820_n N_VGND_c_949_n 0.0116628f $X=5.775 $Y=0.615 $X2=0
+ $Y2=0
cc_516 N_A_27_82#_c_821_n N_VGND_c_949_n 0.0115161f $X=6.64 $Y=0.475 $X2=0 $Y2=0
cc_517 N_A_27_82#_c_822_n N_VGND_c_949_n 0.0499807f $X=7.335 $Y=0.57 $X2=0 $Y2=0
cc_518 N_A_27_82#_c_815_n N_VGND_c_953_n 0.00645633f $X=4.24 $Y=0.555 $X2=0
+ $Y2=0
cc_519 N_A_27_82#_c_857_n N_VGND_c_953_n 0.00322865f $X=5.445 $Y=0.615 $X2=0
+ $Y2=0
cc_520 N_A_27_82#_c_815_n N_VGND_c_954_n 0.00118994f $X=4.24 $Y=0.555 $X2=0
+ $Y2=0
cc_521 N_A_27_82#_c_857_n N_VGND_c_954_n 0.0518121f $X=5.445 $Y=0.615 $X2=0
+ $Y2=0
cc_522 N_A_27_82#_c_820_n N_VGND_c_954_n 0.00471823f $X=5.775 $Y=0.615 $X2=0
+ $Y2=0
cc_523 N_A_27_82#_c_855_n N_VGND_c_955_n 0.0252319f $X=6.475 $Y=0.665 $X2=0
+ $Y2=0
cc_524 N_A_27_82#_c_820_n N_VGND_c_955_n 0.00145033f $X=5.775 $Y=0.615 $X2=0
+ $Y2=0
cc_525 N_A_27_82#_c_821_n N_VGND_c_955_n 0.00151963f $X=6.64 $Y=0.475 $X2=0
+ $Y2=0
