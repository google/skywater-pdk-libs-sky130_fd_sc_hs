* NGSPICE file created from sky130_fd_sc_hs__a21oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_280_107# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=6.5505e+11p pd=6.27e+06u as=4.033e+11p ps=4.05e+06u
M1001 a_131_368# A2 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=1.288e+12p pd=1.126e+07u as=7.392e+11p ps=5.8e+06u
M1002 a_280_107# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.83425e+11p ps=4.82e+06u
M1003 VPWR A1 a_131_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A2 a_280_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_131_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A1 a_280_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_131_368# VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1008 a_131_368# B1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_131_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

