* File: sky130_fd_sc_hs__fahcon_1.pex.spice
* Created: Thu Aug 27 20:46:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A 1 3 4 6 7
c34 7 0 1.4324e-19 $X=0.72 $Y=1.665
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.515 $X2=0.54 $Y2=1.515
r36 7 11 4.82418 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.54 $Y2=1.565
r37 4 10 52.2586 $w=2.99e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.545 $Y=1.765
+ $X2=0.54 $Y2=1.515
r38 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.545 $Y=1.765
+ $X2=0.545 $Y2=2.4
r39 1 10 38.5562 $w=2.99e-07 $l=1.86145e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.54 $Y2=1.515
r40 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.35 $X2=0.495
+ $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_27_100# 1 2 3 4 13 15 16 18 21 27 29 33
+ 37 38 39 44 46 47 48 50 51 54 55 57
c123 57 0 2.01518e-20 $X=1.13 $Y=1.557
c124 33 0 7.413e-20 $X=1.08 $Y=1.515
c125 13 0 1.4324e-19 $X=1.13 $Y=1.765
r126 57 58 31.5515 $w=3.59e-07 $l=2.35e-07 $layer=POLY_cond $X=1.13 $Y=1.557
+ $X2=1.365 $Y2=1.557
r127 54 55 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.81
+ $X2=2.61 $Y2=0.725
r128 50 51 5.26587 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.587 $Y=1.97
+ $X2=2.587 $Y2=1.805
r129 46 47 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=2.115
+ $X2=0.285 $Y2=1.95
r130 42 54 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.61 $Y=0.89 $X2=2.61
+ $Y2=0.81
r131 42 51 31.9541 $w=3.28e-07 $l=9.15e-07 $layer=LI1_cond $X=2.61 $Y=0.89
+ $X2=2.61 $Y2=1.805
r132 40 55 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.53 $Y=0.425
+ $X2=2.53 $Y2=0.725
r133 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=0.34
+ $X2=2.53 $Y2=0.425
r134 38 39 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=2.445 $Y=0.34
+ $X2=1.245 $Y2=0.34
r135 37 48 5.44924 $w=1.87e-07 $l=1.85e-07 $layer=LI1_cond $X=1.16 $Y=0.98
+ $X2=0.975 $Y2=0.98
r136 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.16 $Y=0.425
+ $X2=1.245 $Y2=0.34
r137 36 37 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.16 $Y=0.425
+ $X2=1.16 $Y2=0.98
r138 34 57 6.71309 $w=3.59e-07 $l=5e-08 $layer=POLY_cond $X=1.08 $Y=1.557
+ $X2=1.13 $Y2=1.557
r139 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.515 $X2=1.08 $Y2=1.515
r140 31 48 5.44924 $w=1.87e-07 $l=2.45764e-07 $layer=LI1_cond $X=1.077 $Y=1.18
+ $X2=0.975 $Y2=0.98
r141 31 33 18.1242 $w=2.03e-07 $l=3.35e-07 $layer=LI1_cond $X=1.077 $Y=1.18
+ $X2=1.077 $Y2=1.515
r142 30 44 1.76993 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.08
+ $X2=0.225 $Y2=1.08
r143 29 48 1.11122 $w=2e-07 $l=1e-07 $layer=LI1_cond $X=0.975 $Y=1.08 $X2=0.975
+ $Y2=0.98
r144 29 30 33.8273 $w=1.98e-07 $l=6.1e-07 $layer=LI1_cond $X=0.975 $Y=1.08
+ $X2=0.365 $Y2=1.08
r145 25 46 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=0.285 $Y=2.15
+ $X2=0.285 $Y2=2.115
r146 25 27 19.1594 $w=3.98e-07 $l=6.65e-07 $layer=LI1_cond $X=0.285 $Y=2.15
+ $X2=0.285 $Y2=2.815
r147 23 44 4.67858 $w=2.25e-07 $l=1.24499e-07 $layer=LI1_cond $X=0.17 $Y=1.18
+ $X2=0.225 $Y2=1.08
r148 23 47 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.17 $Y=1.18
+ $X2=0.17 $Y2=1.95
r149 19 44 4.67858 $w=2.25e-07 $l=1e-07 $layer=LI1_cond $X=0.225 $Y=0.98
+ $X2=0.225 $Y2=1.08
r150 19 21 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.225 $Y=0.98
+ $X2=0.225 $Y2=0.645
r151 16 58 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.365 $Y=1.35
+ $X2=1.365 $Y2=1.557
r152 16 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.365 $Y=1.35
+ $X2=1.365 $Y2=0.92
r153 13 57 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.13 $Y=1.765
+ $X2=1.13 $Y2=1.557
r154 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.13 $Y=1.765
+ $X2=1.13 $Y2=2.34
r155 4 50 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=1.825 $X2=2.565 $Y2=1.97
r156 3 46 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.115
r157 3 27 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.815
r158 2 54 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=2.46
+ $Y=0.665 $X2=2.61 $Y2=0.81
r159 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.5 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_336_263# 1 2 8 9 11 15 16 17 18 20 22 24
+ 26 27 33 39 46 47
c116 47 0 2.05468e-19 $X=4.207 $Y=1.805
c117 39 0 1.41326e-19 $X=3.115 $Y=0.405
c118 26 0 7.413e-20 $X=1.775 $Y=1.465
c119 16 0 3.57245e-21 $X=2.75 $Y=0.22
r120 46 47 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=4.207 $Y=1.97
+ $X2=4.207 $Y2=1.805
r121 44 47 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.125 $Y=1.01
+ $X2=4.125 $Y2=1.805
r122 43 44 16.4522 $w=6.93e-07 $l=4.95e-07 $layer=LI1_cond $X=4.387 $Y=0.515
+ $X2=4.387 $Y2=1.01
r123 37 51 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.932 $Y=0.39
+ $X2=2.932 $Y2=0.555
r124 36 39 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=0.405
+ $X2=3.115 $Y2=0.405
r125 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=0.39 $X2=2.95 $Y2=0.39
r126 31 46 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=4.207 $Y=1.972
+ $X2=4.207 $Y2=1.97
r127 31 33 28.4843 $w=3.33e-07 $l=8.28e-07 $layer=LI1_cond $X=4.207 $Y=1.972
+ $X2=4.207 $Y2=2.8
r128 27 43 3.01171 $w=6.93e-07 $l=1.75e-07 $layer=LI1_cond $X=4.387 $Y=0.34
+ $X2=4.387 $Y2=0.515
r129 27 39 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.04 $Y=0.34
+ $X2=3.115 $Y2=0.34
r130 25 26 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.775 $Y=1.315
+ $X2=1.775 $Y2=1.465
r131 24 51 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.825 $Y=0.985
+ $X2=2.825 $Y2=0.555
r132 22 24 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.825 $Y=1.38
+ $X2=2.825 $Y2=0.985
r133 18 22 94.8617 $w=1.88e-07 $l=3.87105e-07 $layer=POLY_cond $X=2.79 $Y=1.75
+ $X2=2.825 $Y2=1.38
r134 18 20 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.79 $Y=1.75
+ $X2=2.79 $Y2=2.245
r135 16 37 26.8759 $w=3.65e-07 $l=1.7e-07 $layer=POLY_cond $X=2.932 $Y=0.22
+ $X2=2.932 $Y2=0.39
r136 16 17 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.75 $Y=0.22
+ $X2=1.87 $Y2=0.22
r137 15 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.795 $Y=0.92
+ $X2=1.795 $Y2=1.315
r138 12 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.795 $Y=0.295
+ $X2=1.87 $Y2=0.22
r139 12 15 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.795 $Y=0.295
+ $X2=1.795 $Y2=0.92
r140 9 11 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.77 $Y=1.75
+ $X2=1.77 $Y2=2.245
r141 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.77 $Y=1.66 $X2=1.77
+ $Y2=1.75
r142 8 26 75.7984 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=1.77 $Y=1.66
+ $X2=1.77 $Y2=1.465
r143 2 46 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.825 $X2=4.21 $Y2=1.97
r144 2 33 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.825 $X2=4.21 $Y2=2.8
r145 1 43 60.6667 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=3
+ $X=4.105 $Y=0.37 $X2=4.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%B 1 2 6 7 9 11 12 13 14 18 21 23 26 27 28
+ 29 31 32 34 36 38 39 41 44 47 48 49 51 56 57
c156 56 0 3.00527e-20 $X=4.9 $Y=1.385
c157 29 0 2.75614e-19 $X=4.435 $Y=1.75
c158 21 0 2.22531e-19 $X=3.43 $Y=0.985
c159 9 0 1.79307e-20 $X=2.385 $Y=0.985
c160 7 0 1.08015e-19 $X=2.385 $Y=1.465
c161 6 0 1.30198e-20 $X=2.34 $Y=2.245
r162 55 57 25.6578 $w=2.63e-07 $l=1.4e-07 $layer=POLY_cond $X=4.9 $Y=1.385
+ $X2=5.04 $Y2=1.385
r163 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.385 $X2=4.9 $Y2=1.385
r164 53 55 16.4943 $w=2.63e-07 $l=9e-08 $layer=POLY_cond $X=4.81 $Y=1.385
+ $X2=4.9 $Y2=1.385
r165 51 56 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.56 $Y=1.365 $X2=4.9
+ $Y2=1.365
r166 46 47 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=3.407 $Y=1.6
+ $X2=3.407 $Y2=1.75
r167 42 57 44.9011 $w=2.63e-07 $l=3.16938e-07 $layer=POLY_cond $X=5.285 $Y=1.22
+ $X2=5.04 $Y2=1.385
r168 42 44 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.285 $Y=1.22
+ $X2=5.285 $Y2=0.69
r169 39 41 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.04 $Y=1.87
+ $X2=5.04 $Y2=2.445
r170 38 39 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.04 $Y=1.78 $X2=5.04
+ $Y2=1.87
r171 37 57 11.6845 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.04 $Y=1.55
+ $X2=5.04 $Y2=1.385
r172 37 38 89.4032 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=5.04 $Y=1.55
+ $X2=5.04 $Y2=1.78
r173 34 53 15.8942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=1.22
+ $X2=4.81 $Y2=1.385
r174 34 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.81 $Y=1.22
+ $X2=4.81 $Y2=0.74
r175 33 49 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.525 $Y=1.475
+ $X2=4.435 $Y2=1.475
r176 32 53 22.5691 $w=2.63e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.735 $Y=1.475
+ $X2=4.81 $Y2=1.385
r177 32 33 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.735 $Y=1.475
+ $X2=4.525 $Y2=1.475
r178 29 49 109.045 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=4.435 $Y=1.75
+ $X2=4.435 $Y2=1.475
r179 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.435 $Y=1.75
+ $X2=4.435 $Y2=2.385
r180 27 49 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.345 $Y=1.475
+ $X2=4.435 $Y2=1.475
r181 27 28 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=4.345 $Y=1.475
+ $X2=3.99 $Y2=1.475
r182 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.915 $Y=1.55
+ $X2=3.99 $Y2=1.475
r183 25 26 761.457 $w=1.5e-07 $l=1.485e-06 $layer=POLY_cond $X=3.915 $Y=1.55
+ $X2=3.915 $Y2=3.035
r184 24 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.49 $Y=3.11 $X2=3.4
+ $Y2=3.11
r185 23 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=3.11
+ $X2=3.915 $Y2=3.035
r186 23 24 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.84 $Y=3.11
+ $X2=3.49 $Y2=3.11
r187 21 46 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.43 $Y=0.985
+ $X2=3.43 $Y2=1.6
r188 18 47 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.4 $Y=2.245
+ $X2=3.4 $Y2=1.75
r189 16 18 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.4 $Y=2.74
+ $X2=3.4 $Y2=2.245
r190 14 48 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.4 $Y=3.035 $X2=3.4
+ $Y2=3.11
r191 13 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.4 $Y=2.83 $X2=3.4
+ $Y2=2.74
r192 13 14 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.4 $Y=2.83
+ $X2=3.4 $Y2=3.035
r193 11 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.31 $Y=3.11 $X2=3.4
+ $Y2=3.11
r194 11 12 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.31 $Y=3.11
+ $X2=2.43 $Y2=3.11
r195 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.385 $Y=1.465
+ $X2=2.385 $Y2=0.985
r196 4 6 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.34 $Y=2.74
+ $X2=2.34 $Y2=2.245
r197 3 7 70.4462 $w=1.95e-07 $l=3.06676e-07 $layer=POLY_cond $X=2.34 $Y=1.75
+ $X2=2.385 $Y2=1.465
r198 3 6 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.34 $Y=1.75
+ $X2=2.34 $Y2=2.245
r199 2 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.34 $Y=3.035
+ $X2=2.43 $Y2=3.11
r200 1 4 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.34 $Y=2.83 $X2=2.34
+ $Y2=2.74
r201 1 2 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.34 $Y=2.83
+ $X2=2.34 $Y2=3.035
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_374_120# 1 2 7 9 12 15 17 19 21 23 24 26
+ 29 32 34 35 41 44 46 48 53 55 57 58 59 60 61 62 69 72 74 82 92
c251 61 0 1.54021e-19 $X=9.215 $Y=0.925
c252 59 0 1.05698e-19 $X=6.815 $Y=0.925
c253 57 0 1.11588e-19 $X=5.855 $Y=0.925
c254 53 0 8.9203e-20 $X=9.58 $Y=1.425
c255 48 0 3.00527e-20 $X=5.702 $Y=1.475
c256 41 0 2.01518e-20 $X=2.01 $Y=1.745
c257 32 0 1.54205e-19 $X=6.977 $Y=1.287
c258 17 0 1.67691e-19 $X=9.5 $Y=1.765
c259 15 0 9.08104e-20 $X=9.455 $Y=0.79
r260 75 92 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=9.36 $Y=0.925
+ $X2=9.56 $Y2=0.925
r261 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0.925
+ $X2=9.36 $Y2=0.925
r262 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0.925
+ $X2=6.96 $Y2=0.925
r263 69 86 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6 $Y=0.925 $X2=5.75
+ $Y2=0.925
r264 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0.925 $X2=6
+ $Y2=0.925
r265 64 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.925
r266 62 71 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=0.925
+ $X2=6.96 $Y2=0.925
r267 61 74 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=0.925
+ $X2=9.36 $Y2=0.925
r268 61 62 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=9.215 $Y=0.925
+ $X2=7.105 $Y2=0.925
r269 60 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=0.925
+ $X2=6 $Y2=0.925
r270 59 71 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=0.925
+ $X2=6.96 $Y2=0.925
r271 59 60 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=6.815 $Y=0.925
+ $X2=6.145 $Y2=0.925
r272 58 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=0.925
+ $X2=2.16 $Y2=0.925
r273 57 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.855 $Y=0.925
+ $X2=6 $Y2=0.925
r274 57 58 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=5.855 $Y=0.925
+ $X2=2.305 $Y2=0.925
r275 53 55 9.38152 $w=2.13e-07 $l=1.65e-07 $layer=LI1_cond $X=9.582 $Y=1.425
+ $X2=9.582 $Y2=1.26
r276 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.58
+ $Y=1.425 $X2=9.58 $Y2=1.425
r277 51 72 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=6.947 $Y=1.13
+ $X2=6.947 $Y2=0.925
r278 46 48 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.702 $Y=1.64
+ $X2=5.702 $Y2=1.475
r279 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.735
+ $Y=1.64 $X2=5.735 $Y2=1.64
r280 43 82 12.8415 $w=3.48e-07 $l=3.9e-07 $layer=LI1_cond $X=2.1 $Y=1.15 $X2=2.1
+ $Y2=0.76
r281 43 44 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=2.1 $Y=1.15
+ $X2=2.1 $Y2=1.325
r282 39 41 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.775 $Y=1.745
+ $X2=2.01 $Y2=1.745
r283 37 92 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.56 $Y=1.04
+ $X2=9.56 $Y2=0.925
r284 37 55 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.56 $Y=1.04
+ $X2=9.56 $Y2=1.26
r285 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.985
+ $Y=1.295 $X2=6.985 $Y2=1.295
r286 32 51 6.1958 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=6.977 $Y=1.287
+ $X2=6.977 $Y2=1.13
r287 32 34 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=6.977 $Y=1.287
+ $X2=6.977 $Y2=1.295
r288 30 86 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.75 $Y=1.04
+ $X2=5.75 $Y2=0.925
r289 30 48 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.75 $Y=1.04
+ $X2=5.75 $Y2=1.475
r290 29 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=1.66
+ $X2=2.01 $Y2=1.745
r291 29 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.01 $Y=1.66
+ $X2=2.01 $Y2=1.325
r292 24 26 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=1.86 $Y=2.65
+ $X2=3.095 $Y2=2.65
r293 23 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.775 $Y=2.565
+ $X2=1.86 $Y2=2.65
r294 22 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=1.83
+ $X2=1.775 $Y2=1.745
r295 22 23 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.775 $Y=1.83
+ $X2=1.775 $Y2=2.565
r296 21 35 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.985 $Y=1.13
+ $X2=6.985 $Y2=1.295
r297 17 54 66.6686 $w=3e-07 $l=3.69703e-07 $layer=POLY_cond $X=9.5 $Y=1.765
+ $X2=9.562 $Y2=1.425
r298 17 19 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.5 $Y=1.765
+ $X2=9.5 $Y2=2.26
r299 13 54 38.5519 $w=3e-07 $l=2.11849e-07 $layer=POLY_cond $X=9.455 $Y=1.26
+ $X2=9.562 $Y2=1.425
r300 13 15 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=9.455 $Y=1.26 $X2=9.455
+ $Y2=0.79
r301 12 21 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.925 $Y=0.69
+ $X2=6.925 $Y2=1.13
r302 7 47 75.7395 $w=2.92e-07 $l=4.44668e-07 $layer=POLY_cond $X=5.575 $Y=2.03
+ $X2=5.692 $Y2=1.64
r303 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.575 $Y=2.03
+ $X2=5.575 $Y2=2.525
r304 2 26 600 $w=1.7e-07 $l=9.32939e-07 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=1.825 $X2=3.095 $Y2=2.65
r305 1 82 91 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.6 $X2=2.09 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_369_365# 1 2 9 11 13 16 18 20 22 23 25 28
+ 33 34 35 36 43 45 52 53 58
c168 53 0 6.54889e-20 $X=8.64 $Y=1.465
c169 52 0 1.54021e-19 $X=8.64 $Y=1.465
c170 28 0 1.30198e-20 $X=2.115 $Y=2.195
c171 23 0 8.9203e-20 $X=9.05 $Y=1.555
c172 9 0 1.54205e-19 $X=6.215 $Y=0.69
r173 52 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.64 $Y=1.465
+ $X2=8.64 $Y2=1.555
r174 52 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.64 $Y=1.465
+ $X2=8.64 $Y2=1.3
r175 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.64
+ $Y=1.465 $X2=8.64 $Y2=1.465
r176 46 53 7.95652 $w=3.68e-07 $l=2.95973e-07 $layer=LI1_cond $X=8.88 $Y=1.665
+ $X2=8.64 $Y2=1.54
r177 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.665
r178 43 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.445
+ $Y=1.715 $X2=6.445 $Y2=1.715
r179 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r180 39 58 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.11 $Y=1.665
+ $X2=3.11 $Y2=0.81
r181 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r182 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=1.665
+ $X2=6.48 $Y2=1.665
r183 35 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=8.88 $Y2=1.665
r184 35 36 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=6.625 $Y2=1.665
r185 34 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r186 33 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=6.48 $Y2=1.665
r187 33 34 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=3.265 $Y2=1.665
r188 32 39 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.11 $Y=2.225
+ $X2=3.11 $Y2=1.665
r189 28 30 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.115 $Y=2.195
+ $X2=2.115 $Y2=2.31
r190 26 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.31
+ $X2=2.115 $Y2=2.31
r191 25 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.945 $Y=2.31
+ $X2=3.11 $Y2=2.225
r192 25 26 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.945 $Y=2.31
+ $X2=2.2 $Y2=2.31
r193 20 23 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=9.05 $Y=1.765
+ $X2=9.05 $Y2=1.555
r194 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.05 $Y=1.765
+ $X2=9.05 $Y2=2.26
r195 19 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.805 $Y=1.555
+ $X2=8.64 $Y2=1.555
r196 18 23 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.96 $Y=1.555 $X2=9.05
+ $Y2=1.555
r197 18 19 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=8.96 $Y=1.555
+ $X2=8.805 $Y2=1.555
r198 16 54 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=8.645 $Y=0.79
+ $X2=8.645 $Y2=1.3
r199 11 49 58.2777 $w=3.79e-07 $l=3.80657e-07 $layer=POLY_cond $X=6.23 $Y=2.03
+ $X2=6.375 $Y2=1.715
r200 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.23 $Y=2.03
+ $X2=6.23 $Y2=2.525
r201 7 49 39.2012 $w=3.79e-07 $l=2.31571e-07 $layer=POLY_cond $X=6.215 $Y=1.55
+ $X2=6.375 $Y2=1.715
r202 7 9 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.215 $Y=1.55
+ $X2=6.215 $Y2=0.69
r203 2 28 600 $w=1.7e-07 $l=4.86621e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.825 $X2=2.115 $Y2=2.195
r204 1 58 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.9
+ $Y=0.665 $X2=3.11 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%CI 5 8 10 12 13 15 16 17 18 25
c65 25 0 6.54889e-20 $X=7.955 $Y=1.492
c66 8 0 2.79202e-20 $X=7.625 $Y=0.69
r67 23 25 19.0481 $w=2.91e-07 $l=1.15e-07 $layer=POLY_cond $X=7.84 $Y=1.492
+ $X2=7.955 $Y2=1.492
r68 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.84
+ $Y=1.385 $X2=7.84 $Y2=1.385
r69 21 23 35.6117 $w=2.91e-07 $l=2.15e-07 $layer=POLY_cond $X=7.625 $Y=1.492
+ $X2=7.84 $Y2=1.492
r70 18 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.84 $Y=1.295 $X2=7.84
+ $Y2=1.385
r71 16 17 41.3838 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=7.442 $Y=1.79
+ $X2=7.442 $Y2=1.885
r72 13 25 29.8144 $w=2.91e-07 $l=3.50634e-07 $layer=POLY_cond $X=8.135 $Y=1.22
+ $X2=7.955 $Y2=1.492
r73 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.135 $Y=1.22
+ $X2=8.135 $Y2=0.74
r74 10 25 18.2534 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=7.955 $Y=1.765
+ $X2=7.955 $Y2=1.492
r75 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.955 $Y=1.765
+ $X2=7.955 $Y2=2.4
r76 6 21 18.2534 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=7.625 $Y=1.22
+ $X2=7.625 $Y2=1.492
r77 6 8 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.625 $Y=1.22
+ $X2=7.625 $Y2=0.69
r78 5 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.45 $Y=2.46
+ $X2=7.45 $Y2=1.885
r79 1 21 31.4708 $w=2.91e-07 $l=1.9e-07 $layer=POLY_cond $X=7.435 $Y=1.492
+ $X2=7.625 $Y2=1.492
r80 1 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.435 $Y=1.55
+ $X2=7.435 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_1606_368# 1 2 3 12 15 16 18 20 22 25 29
+ 33 36 39 40 42 45 46 50 51
c122 40 0 1.25754e-19 $X=8.18 $Y=2.405
c123 39 0 2.79202e-20 $X=8.18 $Y=1.82
r124 51 53 0.995868 $w=2.42e-07 $l=5e-09 $layer=POLY_cond $X=10.12 $Y=1.425
+ $X2=10.115 $Y2=1.425
r125 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.12
+ $Y=1.425 $X2=10.12 $Y2=1.425
r126 47 50 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=9.945 $Y=1.425
+ $X2=10.12 $Y2=1.425
r127 45 46 9.33757 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.795 $Y=1.985
+ $X2=9.795 $Y2=1.82
r128 42 43 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=8.345 $Y=0.965
+ $X2=8.345 $Y2=1.13
r129 39 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.26 $Y=1.82
+ $X2=8.26 $Y2=1.13
r130 37 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.945 $Y=1.59
+ $X2=9.945 $Y2=1.425
r131 37 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.945 $Y=1.59
+ $X2=9.945 $Y2=1.82
r132 35 45 1.78139 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=9.795 $Y=2.055
+ $X2=9.795 $Y2=1.985
r133 35 36 6.74385 $w=4.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.795 $Y=2.055
+ $X2=9.795 $Y2=2.32
r134 34 40 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.345 $Y=2.405
+ $X2=8.18 $Y2=2.405
r135 33 36 8.97637 $w=1.7e-07 $l=2.74226e-07 $layer=LI1_cond $X=9.56 $Y=2.405
+ $X2=9.795 $Y2=2.32
r136 33 34 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=9.56 $Y=2.405
+ $X2=8.345 $Y2=2.405
r137 27 42 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=8.345 $Y=0.96
+ $X2=8.345 $Y2=0.965
r138 27 29 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=8.345 $Y=0.96
+ $X2=8.345 $Y2=0.515
r139 23 40 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.18 $Y=2.49
+ $X2=8.18 $Y2=2.405
r140 23 25 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.18 $Y=2.49
+ $X2=8.18 $Y2=2.815
r141 22 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.18 $Y=1.985
+ $X2=8.18 $Y2=1.82
r142 20 40 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.18 $Y=2.32
+ $X2=8.18 $Y2=2.405
r143 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.18 $Y=2.32
+ $X2=8.18 $Y2=1.985
r144 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=10.51 $Y=1.885
+ $X2=10.51 $Y2=2.46
r145 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.51 $Y=1.795
+ $X2=10.51 $Y2=1.885
r146 14 51 77.6777 $w=2.42e-07 $l=4.65242e-07 $layer=POLY_cond $X=10.51 $Y=1.59
+ $X2=10.12 $Y2=1.425
r147 14 15 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=10.51 $Y=1.59
+ $X2=10.51 $Y2=1.795
r148 10 53 13.9682 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.115 $Y=1.26
+ $X2=10.115 $Y2=1.425
r149 10 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=10.115 $Y=1.26
+ $X2=10.115 $Y2=0.79
r150 3 45 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.575
+ $Y=1.84 $X2=9.725 $Y2=1.985
r151 2 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.03
+ $Y=1.84 $X2=8.18 $Y2=2.815
r152 2 22 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.03
+ $Y=1.84 $X2=8.18 $Y2=1.985
r153 1 42 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.21
+ $Y=0.37 $X2=8.35 $Y2=0.965
r154 1 29 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.21
+ $Y=0.37 $X2=8.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_1744_94# 1 2 7 9 12 15 17 18 19 23 24 25
+ 31 32 35 37
c104 25 0 9.08104e-20 $X=10.325 $Y=0.665
r105 35 37 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=10.952 $Y=1.465
+ $X2=10.952 $Y2=1.3
r106 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.975
+ $Y=1.465 $X2=10.975 $Y2=1.465
r107 31 32 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=9.247 $Y=1.985
+ $X2=9.247 $Y2=1.82
r108 26 37 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=10.895 $Y=0.75
+ $X2=10.895 $Y2=1.3
r109 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.81 $Y=0.665
+ $X2=10.895 $Y2=0.75
r110 24 25 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=10.81 $Y=0.665
+ $X2=10.325 $Y2=0.665
r111 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.24 $Y=0.58
+ $X2=10.325 $Y2=0.665
r112 22 23 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.24 $Y=0.425
+ $X2=10.24 $Y2=0.58
r113 20 32 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=9.22 $Y=1.38
+ $X2=9.22 $Y2=1.82
r114 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.155 $Y=0.34
+ $X2=10.24 $Y2=0.425
r115 18 19 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=10.155 $Y=0.34
+ $X2=9.105 $Y2=0.34
r116 15 20 13.83 $w=2.47e-07 $l=3.69648e-07 $layer=LI1_cond $X=8.94 $Y=1.172
+ $X2=9.22 $Y2=1.38
r117 15 17 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.94 $Y=0.965
+ $X2=8.94 $Y2=0.615
r118 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.94 $Y=0.425
+ $X2=9.105 $Y2=0.34
r119 14 17 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=8.94 $Y=0.425
+ $X2=8.94 $Y2=0.615
r120 10 36 38.6549 $w=2.86e-07 $l=1.88348e-07 $layer=POLY_cond $X=11.025 $Y=1.3
+ $X2=10.975 $Y2=1.465
r121 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.025 $Y=1.3
+ $X2=11.025 $Y2=0.74
r122 7 36 61.4066 $w=2.86e-07 $l=3.19374e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=10.975 $Y2=1.465
r123 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=11.015 $Y2=2.4
r124 2 31 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.125
+ $Y=1.84 $X2=9.275 $Y2=1.985
r125 1 17 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.47 $X2=8.94 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%VPWR 1 2 3 4 17 23 29 35 38 39 40 42 54 63
+ 64 67 70 73
r95 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r96 70 71 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 64 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r99 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r100 61 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.9 $Y=3.33
+ $X2=10.775 $Y2=3.33
r101 61 63 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.9 $Y=3.33
+ $X2=11.28 $Y2=3.33
r102 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r103 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r104 57 60 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r105 56 59 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r106 56 57 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r107 54 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=10.775 $Y2=3.33
r108 54 59 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=10.32 $Y2=3.33
r109 53 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r110 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r111 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 49 52 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r114 47 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=4.71 $Y2=3.33
r115 47 49 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 46 71 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 46 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 45 46 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r120 43 45 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r121 42 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.71 $Y2=3.33
r122 42 45 218.23 $w=1.68e-07 $l=3.345e-06 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 40 53 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=7.44 $Y2=3.33
r124 40 50 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 38 52 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.645 $Y=3.33
+ $X2=7.44 $Y2=3.33
r126 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.645 $Y=3.33
+ $X2=7.73 $Y2=3.33
r127 37 56 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.815 $Y=3.33
+ $X2=7.92 $Y2=3.33
r128 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=3.33
+ $X2=7.73 $Y2=3.33
r129 33 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.775 $Y=3.245
+ $X2=10.775 $Y2=3.33
r130 33 35 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=10.775 $Y=3.245
+ $X2=10.775 $Y2=2.265
r131 29 32 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.73 $Y=2.105
+ $X2=7.73 $Y2=2.815
r132 27 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.73 $Y=3.245
+ $X2=7.73 $Y2=3.33
r133 27 32 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.73 $Y=3.245
+ $X2=7.73 $Y2=2.815
r134 23 26 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.71 $Y=1.97
+ $X2=4.71 $Y2=2.385
r135 21 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.71 $Y=3.245
+ $X2=4.71 $Y2=3.33
r136 21 26 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.71 $Y=3.245
+ $X2=4.71 $Y2=2.385
r137 17 20 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.82 $Y=2.115
+ $X2=0.82 $Y2=2.815
r138 15 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=3.33
r139 15 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.815
r140 4 35 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=10.585
+ $Y=1.96 $X2=10.735 $Y2=2.265
r141 3 32 400 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=7.525
+ $Y=1.96 $X2=7.73 $Y2=2.815
r142 3 29 400 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=7.525
+ $Y=1.96 $X2=7.73 $Y2=2.105
r143 2 26 300 $w=1.7e-07 $l=6.5238e-07 $layer=licon1_PDIFF $count=2 $X=4.51
+ $Y=1.825 $X2=4.71 $Y2=2.385
r144 2 23 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.825 $X2=4.71 $Y2=1.97
r145 1 20 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.84 $X2=0.82 $Y2=2.815
r146 1 17 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=0.62
+ $Y=1.84 $X2=0.82 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_241_368# 1 2 3 4 16 18 23 25 26 29 33 35
c72 25 0 1.69282e-19 $X=3.46 $Y=2.99
r73 34 35 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.547 $Y=1.32
+ $X2=1.547 $Y2=1.49
r74 33 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.435 $Y=1.85
+ $X2=1.435 $Y2=1.49
r75 29 32 38.1953 $w=3.48e-07 $l=1.16e-06 $layer=LI1_cond $X=3.635 $Y=0.81
+ $X2=3.635 $Y2=1.97
r76 27 32 30.7867 $w=3.48e-07 $l=9.35e-07 $layer=LI1_cond $X=3.635 $Y=2.905
+ $X2=3.635 $Y2=1.97
r77 25 27 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=3.46 $Y=2.99
+ $X2=3.635 $Y2=2.905
r78 25 26 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=3.46 $Y=2.99
+ $X2=1.52 $Y2=2.99
r79 23 34 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.58 $Y=0.76
+ $X2=1.58 $Y2=1.32
r80 16 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.015
+ $X2=1.355 $Y2=1.85
r81 16 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.355 $Y=2.015
+ $X2=1.355 $Y2=2.695
r82 14 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.355 $Y=2.905
+ $X2=1.52 $Y2=2.99
r83 14 18 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.355 $Y=2.905
+ $X2=1.355 $Y2=2.695
r84 4 32 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.475
+ $Y=1.825 $X2=3.625 $Y2=1.97
r85 3 18 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.84 $X2=1.355 $Y2=2.695
r86 3 16 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=1.205
+ $Y=1.84 $X2=1.355 $Y2=2.015
r87 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.665 $X2=3.645 $Y2=0.81
r88 1 23 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=1.44
+ $Y=0.6 $X2=1.58 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_1023_389# 1 2 9 14 15 17 20 21 24
c56 17 0 1.05698e-19 $X=5.985 $Y=0.555
r57 22 24 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.315 $Y=1.22
+ $X2=5.41 $Y2=1.22
r58 20 21 7.76373 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.265 $Y=2.12
+ $X2=5.265 $Y2=1.975
r59 15 17 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=5.495 $Y=0.515
+ $X2=5.985 $Y2=0.515
r60 14 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=1.135
+ $X2=5.41 $Y2=1.22
r61 13 15 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.41 $Y=0.64
+ $X2=5.495 $Y2=0.515
r62 13 14 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.41 $Y=0.64
+ $X2=5.41 $Y2=1.135
r63 11 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=1.305
+ $X2=5.315 $Y2=1.22
r64 11 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.315 $Y=1.305
+ $X2=5.315 $Y2=1.975
r65 7 20 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=5.265 $Y=2.14 $X2=5.265
+ $Y2=2.12
r66 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.265 $Y=2.14
+ $X2=5.265 $Y2=2.46
r67 2 20 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=5.115
+ $Y=1.945 $X2=5.265 $Y2=2.12
r68 2 9 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=5.115
+ $Y=1.945 $X2=5.265 $Y2=2.46
r69 1 17 91 $w=1.7e-07 $l=7.11512e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.37 $X2=5.985 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%COUT_N 1 2 12 13 18 20
r52 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.485 $Y=1.21
+ $X2=6.485 $Y2=0.515
r53 15 18 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.09 $Y=1.295
+ $X2=6.485 $Y2=1.295
r54 12 13 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.982 $Y=2.25
+ $X2=5.982 $Y2=2.085
r55 9 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=1.38 $X2=6.09
+ $Y2=1.295
r56 9 13 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.09 $Y=1.38
+ $X2=6.09 $Y2=2.085
r57 2 12 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=5.65
+ $Y=2.105 $X2=5.955 $Y2=2.25
r58 1 20 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=6.29
+ $Y=0.37 $X2=6.485 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_1261_421# 1 2 7 15 18 19
r47 18 19 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=7.39 $Y=2.085
+ $X2=7.39 $Y2=0.96
r48 13 19 7.30505 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=0.795
+ $X2=7.41 $Y2=0.96
r49 13 15 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.41 $Y=0.795
+ $X2=7.41 $Y2=0.515
r50 9 12 10.6147 $w=8.83e-07 $l=7.7e-07 $layer=LI1_cond $X=6.455 $Y=2.527
+ $X2=7.225 $Y2=2.527
r51 7 18 12.0616 $w=8.85e-07 $l=4.82632e-07 $layer=LI1_cond $X=7.305 $Y=2.527
+ $X2=7.39 $Y2=2.085
r52 7 12 1.10282 $w=8.83e-07 $l=8e-08 $layer=LI1_cond $X=7.305 $Y=2.527
+ $X2=7.225 $Y2=2.527
r53 2 12 200 $w=1.7e-07 $l=9.89848e-07 $layer=licon1_PDIFF $count=3 $X=6.305
+ $Y=2.105 $X2=7.225 $Y2=2.25
r54 2 9 200 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=3 $X=6.305
+ $Y=2.105 $X2=6.455 $Y2=2.25
r55 1 15 91 $w=1.7e-07 $l=4.77022e-07 $layer=licon1_NDIFF $count=2 $X=7 $Y=0.37
+ $X2=7.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%A_1719_368# 1 2 3 10 14 16 17 21 25 27 33
c66 33 0 1.67691e-19 $X=10.54 $Y=1.845
r67 27 29 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.74 $Y=2.825
+ $X2=8.74 $Y2=2.955
r68 25 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.54 $Y=1.76
+ $X2=10.54 $Y2=1.845
r69 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.54 $Y=1.09
+ $X2=10.54 $Y2=1.76
r70 21 23 32.0876 $w=2.53e-07 $l=7.1e-07 $layer=LI1_cond $X=10.327 $Y=2.105
+ $X2=10.327 $Y2=2.815
r71 19 23 2.48566 $w=2.53e-07 $l=5.5e-08 $layer=LI1_cond $X=10.327 $Y=2.87
+ $X2=10.327 $Y2=2.815
r72 18 33 13.8963 $w=1.68e-07 $l=2.13e-07 $layer=LI1_cond $X=10.327 $Y=1.845
+ $X2=10.54 $Y2=1.845
r73 18 21 7.90892 $w=2.53e-07 $l=1.75e-07 $layer=LI1_cond $X=10.327 $Y=1.93
+ $X2=10.327 $Y2=2.105
r74 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.455 $Y=1.005
+ $X2=10.54 $Y2=1.09
r75 16 17 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=10.455 $Y=1.005
+ $X2=9.985 $Y2=1.005
r76 12 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.9 $Y=0.92
+ $X2=9.985 $Y2=1.005
r77 12 14 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=9.9 $Y=0.92 $X2=9.9
+ $Y2=0.84
r78 11 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.905 $Y=2.955
+ $X2=8.74 $Y2=2.955
r79 10 19 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=10.2 $Y=2.955
+ $X2=10.327 $Y2=2.87
r80 10 11 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=10.2 $Y=2.955
+ $X2=8.905 $Y2=2.955
r81 3 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.96 $X2=10.285 $Y2=2.815
r82 3 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.96 $X2=10.285 $Y2=2.105
r83 2 27 600 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=8.595
+ $Y=1.84 $X2=8.74 $Y2=2.825
r84 1 14 182 $w=1.7e-07 $l=5.23259e-07 $layer=licon1_NDIFF $count=1 $X=9.53
+ $Y=0.47 $X2=9.9 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%SUM 1 2 9 13 14 15 16 23 32
r26 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=11.255 $Y=2
+ $X2=11.255 $Y2=2.035
r27 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=11.255 $Y=2.405
+ $X2=11.255 $Y2=2.775
r28 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=2
r29 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=1.82
r30 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.405
r31 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.035
r32 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.35 $Y=1.13
+ $X2=11.35 $Y2=1.82
r33 7 13 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=11.295 $Y=0.99
+ $X2=11.295 $Y2=1.13
r34 7 9 19.5504 $w=2.78e-07 $l=4.75e-07 $layer=LI1_cond $X=11.295 $Y=0.99
+ $X2=11.295 $Y2=0.515
r35 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=1.985
r36 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=2.815
r37 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.1
+ $Y=0.37 $X2=11.24 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCON_1%VGND 1 2 3 4 14 17 21 24 25 29 31 37 44 52
+ 59 60 63 66 70
r108 70 73 9.3636 $w=3.98e-07 $l=3.25e-07 $layer=LI1_cond $X=10.695 $Y=0
+ $X2=10.695 $Y2=0.325
r109 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r110 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r111 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r112 60 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r113 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r114 57 70 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.895 $Y=0 $X2=10.695
+ $Y2=0
r115 57 59 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.28 $Y2=0
r116 56 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r117 56 67 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=7.92 $Y2=0
r118 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r119 53 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=7.87
+ $Y2=0
r120 53 55 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=7.995 $Y=0
+ $X2=10.32 $Y2=0
r121 52 70 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.495 $Y=0 $X2=10.695
+ $Y2=0
r122 52 55 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.32 $Y2=0
r123 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r124 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r125 48 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r126 47 50 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r127 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r128 45 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=5.03
+ $Y2=0
r129 45 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=5.52 $Y2=0
r130 44 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.87
+ $Y2=0
r131 44 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r132 43 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r133 42 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r134 40 43 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.72 $Y=0 $X2=4.56
+ $Y2=0
r135 39 42 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=4.56
+ $Y2=0
r136 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r137 37 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.905 $Y=0 $X2=5.03
+ $Y2=0
r138 37 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.905 $Y=0 $X2=4.56
+ $Y2=0
r139 35 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r140 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r141 31 51 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r142 31 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r143 26 29 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.63 $Y=0.645
+ $X2=0.725 $Y2=0.645
r144 24 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r145 24 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.63
+ $Y2=0
r146 23 39 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.72
+ $Y2=0
r147 23 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.63
+ $Y2=0
r148 19 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0
r149 19 21 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0.495
r150 15 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r151 15 17 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.655
r152 14 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0.48
+ $X2=0.63 $Y2=0.645
r153 13 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.085
+ $X2=0.63 $Y2=0
r154 13 14 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.63 $Y=0.085
+ $X2=0.63 $Y2=0.48
r155 4 73 182 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_NDIFF $count=1 $X=10.19
+ $Y=0.47 $X2=10.695 $Y2=0.325
r156 3 21 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=7.7
+ $Y=0.37 $X2=7.91 $Y2=0.495
r157 2 17 182 $w=1.7e-07 $l=3.65992e-07 $layer=licon1_NDIFF $count=1 $X=4.885
+ $Y=0.37 $X2=5.07 $Y2=0.655
r158 1 29 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.5 $X2=0.725 $Y2=0.645
.ends

