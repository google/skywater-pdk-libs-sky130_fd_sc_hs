* File: sky130_fd_sc_hs__clkbuf_8.spice
* Created: Thu Aug 27 20:35:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__clkbuf_8.pex.spice"
.subckt sky130_fd_sc_hs__clkbuf_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_125_368#_M1007_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.3
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g N_A_125_368#_M1007_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.08295 AS=0.0588 PD=0.815 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75004 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1010_d N_A_125_368#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.08295 AS=0.06405 PD=0.815 PS=0.725 NRD=12.852 NRS=7.14 M=1 R=2.8
+ SA=75001.3 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_125_368#_M1002_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.06405 PD=0.84 PS=0.725 NRD=19.992 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1002_d N_A_125_368#_M1003_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.0588 PD=0.84 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_125_368#_M1004_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.7 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1004_d N_A_125_368#_M1006_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.1 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_125_368#_M1008_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=9.996 NRS=0 M=1 R=2.8 SA=75003.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1008_d N_A_125_368#_M1018_g N_X_M1018_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=9.996 NRS=0 M=1 R=2.8 SA=75004.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_125_368#_M1019_g N_X_M1018_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_A_125_368#_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3808 AS=0.1708 PD=2.92 PS=1.425 NRD=9.6727 NRS=2.6201 M=1 R=7.46667
+ SA=75000.3 SB=75004.4 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g N_A_125_368#_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.224 AS=0.1708 PD=1.52 PS=1.425 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75004 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1016_d N_A_125_368#_M1001_g N_X_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.3 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A_125_368#_M1005_g N_X_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75003 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1005_d N_A_125_368#_M1009_g N_X_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.2 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1012_d N_A_125_368#_M1012_g N_X_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1012_d N_A_125_368#_M1013_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A_125_368#_M1014_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1014_d N_A_125_368#_M1015_g N_X_M1015_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.1764 PD=1.47 PS=1.435 NRD=10.5395 NRS=2.6201 M=1 R=7.46667
+ SA=75004 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1017_d N_A_125_368#_M1017_g N_X_M1015_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.1764 PD=2.83 PS=1.435 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75004.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_hs__clkbuf_8.pxi.spice"
*
.ends
*
*
