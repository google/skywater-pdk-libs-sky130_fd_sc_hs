* File: sky130_fd_sc_hs__o2111a_2.pxi.spice
* Created: Tue Sep  1 20:13:04 2020
* 
x_PM_SKY130_FD_SC_HS__O2111A_2%A1 N_A1_c_73_n N_A1_c_77_n N_A1_M1000_g
+ N_A1_M1010_g A1 A1 N_A1_c_75_n PM_SKY130_FD_SC_HS__O2111A_2%A1
x_PM_SKY130_FD_SC_HS__O2111A_2%A2 N_A2_c_97_n N_A2_M1003_g N_A2_c_98_n
+ N_A2_M1001_g A2 PM_SKY130_FD_SC_HS__O2111A_2%A2
x_PM_SKY130_FD_SC_HS__O2111A_2%B1 N_B1_c_125_n N_B1_M1009_g N_B1_c_126_n
+ N_B1_M1013_g B1 PM_SKY130_FD_SC_HS__O2111A_2%B1
x_PM_SKY130_FD_SC_HS__O2111A_2%C1 N_C1_M1006_g N_C1_c_158_n N_C1_M1007_g C1
+ PM_SKY130_FD_SC_HS__O2111A_2%C1
x_PM_SKY130_FD_SC_HS__O2111A_2%D1 N_D1_M1011_g N_D1_c_197_n N_D1_M1008_g D1
+ N_D1_c_195_n N_D1_c_196_n PM_SKY130_FD_SC_HS__O2111A_2%D1
x_PM_SKY130_FD_SC_HS__O2111A_2%A_236_368# N_A_236_368#_M1011_d
+ N_A_236_368#_M1003_d N_A_236_368#_M1007_d N_A_236_368#_c_240_n
+ N_A_236_368#_M1004_g N_A_236_368#_M1002_g N_A_236_368#_c_241_n
+ N_A_236_368#_M1005_g N_A_236_368#_M1012_g N_A_236_368#_c_242_n
+ N_A_236_368#_c_243_n N_A_236_368#_c_253_n N_A_236_368#_c_244_n
+ N_A_236_368#_c_261_n N_A_236_368#_c_234_n N_A_236_368#_c_235_n
+ N_A_236_368#_c_236_n N_A_236_368#_c_237_n N_A_236_368#_c_238_n
+ N_A_236_368#_c_264_n N_A_236_368#_c_239_n
+ PM_SKY130_FD_SC_HS__O2111A_2%A_236_368#
x_PM_SKY130_FD_SC_HS__O2111A_2%VPWR N_VPWR_M1000_s N_VPWR_M1009_d N_VPWR_M1008_d
+ N_VPWR_M1005_s N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n
+ N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n
+ VPWR N_VPWR_c_348_n N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_338_n
+ PM_SKY130_FD_SC_HS__O2111A_2%VPWR
x_PM_SKY130_FD_SC_HS__O2111A_2%X N_X_M1002_s N_X_M1004_d N_X_c_399_n N_X_c_400_n
+ N_X_c_396_n X X X PM_SKY130_FD_SC_HS__O2111A_2%X
x_PM_SKY130_FD_SC_HS__O2111A_2%A_54_74# N_A_54_74#_M1010_s N_A_54_74#_M1001_d
+ N_A_54_74#_c_427_n N_A_54_74#_c_428_n N_A_54_74#_c_433_n N_A_54_74#_c_439_n
+ N_A_54_74#_c_429_n PM_SKY130_FD_SC_HS__O2111A_2%A_54_74#
x_PM_SKY130_FD_SC_HS__O2111A_2%VGND N_VGND_M1010_d N_VGND_M1002_d N_VGND_M1012_d
+ N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n N_VGND_c_457_n VGND
+ N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n
+ N_VGND_c_463_n PM_SKY130_FD_SC_HS__O2111A_2%VGND
cc_1 VNB N_A1_c_73_n 0.0782236f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.385
cc_2 VNB A1 0.0291142f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A1_c_75_n 0.023452f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.22
cc_4 VNB N_A2_c_97_n 0.0392615f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.385
cc_5 VNB N_A2_c_98_n 0.0186009f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.34
cc_6 VNB A2 0.00596829f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_7 VNB N_B1_c_125_n 0.0378482f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.385
cc_8 VNB N_B1_c_126_n 0.0183068f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.34
cc_9 VNB B1 0.00892781f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_10 VNB N_C1_M1006_g 0.026905f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.765
cc_11 VNB N_C1_c_158_n 0.0282117f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.34
cc_12 VNB C1 0.0121385f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_13 VNB N_D1_M1011_g 0.030729f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.765
cc_14 VNB N_D1_c_195_n 0.0377201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D1_c_196_n 0.00305137f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.22
cc_16 VNB N_A_236_368#_M1002_g 0.0223898f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_17 VNB N_A_236_368#_M1012_g 0.0266858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_236_368#_c_234_n 0.00994708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_236_368#_c_235_n 0.0187701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_236_368#_c_236_n 0.00248805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_236_368#_c_237_n 0.0094184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_236_368#_c_238_n 4.18697e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_236_368#_c_239_n 0.081062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_338_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_396_n 0.00270411f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_26 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_27 VNB X 0.00448002f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_28 VNB N_A_54_74#_c_427_n 0.00716827f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_29 VNB N_A_54_74#_c_428_n 0.0217137f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_A_54_74#_c_429_n 0.00280313f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_31 VNB N_VGND_c_454_n 0.00460613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_455_n 0.0145024f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_33 VNB N_VGND_c_456_n 0.0109665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_457_n 0.0516149f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_35 VNB N_VGND_c_458_n 0.0232895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_459_n 0.0643439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_460_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_461_n 0.00866122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_462_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_463_n 0.308027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A1_c_73_n 0.0100934f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.385
cc_42 VPB N_A1_c_77_n 0.0180428f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.765
cc_43 VPB N_A2_c_97_n 0.0240617f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.385
cc_44 VPB N_B1_c_125_n 0.0250891f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.385
cc_45 VPB N_C1_c_158_n 0.0276421f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=2.34
cc_46 VPB C1 0.00566637f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.74
cc_47 VPB N_D1_c_197_n 0.0175965f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=2.34
cc_48 VPB N_D1_c_195_n 0.0173108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_D1_c_196_n 0.00444844f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.22
cc_50 VPB N_A_236_368#_c_240_n 0.0161702f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_51 VPB N_A_236_368#_c_241_n 0.017345f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_52 VPB N_A_236_368#_c_242_n 0.0100959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_236_368#_c_243_n 0.00357711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_236_368#_c_244_n 0.00359402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_236_368#_c_238_n 0.00340501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_236_368#_c_239_n 0.0169047f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_339_n 0.0613622f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_58 VPB N_VPWR_c_340_n 0.0198828f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_59 VPB N_VPWR_c_341_n 0.018006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_342_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_343_n 0.0693139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_344_n 0.0115308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_345_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_346_n 0.0348258f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_347_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_348_n 0.0220157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_349_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_350_n 0.0155543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_338_n 0.0994504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_X_c_399_n 0.00166049f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_71 VPB N_X_c_400_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_X_c_396_n 8.14144e-19 $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_73 N_A1_c_73_n N_A2_c_97_n 0.0304064f $X=0.595 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_74 N_A1_c_77_n N_A2_c_97_n 0.0532832f $X=0.685 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_75 A1 N_A2_c_97_n 0.00216087f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_76 N_A1_c_75_n N_A2_c_98_n 0.0268292f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_77 N_A1_c_73_n A2 3.68035e-19 $X=0.595 $Y=1.385 $X2=0 $Y2=0
cc_78 A1 A2 0.029889f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A1_c_73_n N_VPWR_c_339_n 0.00704273f $X=0.595 $Y=1.385 $X2=0 $Y2=0
cc_80 N_A1_c_77_n N_VPWR_c_339_n 0.0249128f $X=0.685 $Y=1.765 $X2=0 $Y2=0
cc_81 A1 N_VPWR_c_339_n 0.0196555f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A1_c_77_n N_VPWR_c_346_n 0.00443511f $X=0.685 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A1_c_77_n N_VPWR_c_338_n 0.00460931f $X=0.685 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A1_c_73_n N_A_54_74#_c_427_n 0.00229697f $X=0.595 $Y=1.385 $X2=0 $Y2=0
cc_85 A1 N_A_54_74#_c_427_n 0.0282818f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A1_c_75_n N_A_54_74#_c_428_n 8.37507e-19 $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_87 A1 N_A_54_74#_c_433_n 0.0153343f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A1_c_75_n N_A_54_74#_c_433_n 0.0102656f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_89 N_A1_c_75_n N_VGND_c_454_n 0.0159254f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_90 N_A1_c_75_n N_VGND_c_458_n 0.00383152f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_91 N_A1_c_75_n N_VGND_c_463_n 0.00388149f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_92 N_A2_c_97_n N_B1_c_125_n 0.041652f $X=1.105 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_93 A2 N_B1_c_125_n 4.06701e-19 $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_94 N_A2_c_98_n N_B1_c_126_n 0.0198524f $X=1.27 $Y=1.22 $X2=0 $Y2=0
cc_95 N_A2_c_98_n B1 0.00228667f $X=1.27 $Y=1.22 $X2=0 $Y2=0
cc_96 A2 B1 0.0242365f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A2_c_97_n N_A_236_368#_c_242_n 0.00514342f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_98 A2 N_A_236_368#_c_242_n 0.00356336f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A2_c_97_n N_A_236_368#_c_243_n 0.0108202f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A2_c_97_n N_VPWR_c_339_n 0.00367669f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A2_c_97_n N_VPWR_c_346_n 0.0049405f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A2_c_97_n N_VPWR_c_338_n 0.00508379f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A2_c_97_n N_A_54_74#_c_433_n 9.99496e-19 $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A2_c_98_n N_A_54_74#_c_433_n 0.0126376f $X=1.27 $Y=1.22 $X2=0 $Y2=0
cc_105 A2 N_A_54_74#_c_433_n 0.0228656f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A2_c_98_n N_A_54_74#_c_429_n 0.0026172f $X=1.27 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A2_c_98_n N_VGND_c_454_n 0.0131556f $X=1.27 $Y=1.22 $X2=0 $Y2=0
cc_108 N_A2_c_98_n N_VGND_c_459_n 0.00383152f $X=1.27 $Y=1.22 $X2=0 $Y2=0
cc_109 N_A2_c_98_n N_VGND_c_463_n 0.00384679f $X=1.27 $Y=1.22 $X2=0 $Y2=0
cc_110 N_B1_c_125_n N_C1_M1006_g 0.0179214f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B1_c_126_n N_C1_M1006_g 0.0415061f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_112 B1 N_C1_M1006_g 0.00173356f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B1_c_125_n N_C1_c_158_n 0.0273985f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_114 B1 N_C1_c_158_n 2.54315e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B1_c_125_n C1 0.00366387f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_116 B1 C1 0.0119739f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B1_c_125_n N_A_236_368#_c_242_n 0.00393524f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_118 B1 N_A_236_368#_c_242_n 0.00297112f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B1_c_125_n N_A_236_368#_c_243_n 0.00946384f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_120 N_B1_c_125_n N_A_236_368#_c_253_n 0.0146278f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_121 B1 N_A_236_368#_c_253_n 0.0101041f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B1_c_125_n N_A_236_368#_c_244_n 8.78407e-19 $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_B1_c_125_n N_VPWR_c_340_n 0.00741274f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B1_c_125_n N_VPWR_c_346_n 0.00481995f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B1_c_125_n N_VPWR_c_338_n 0.00508379f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B1_c_125_n N_A_54_74#_c_439_n 6.0983e-19 $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_127 N_B1_c_126_n N_A_54_74#_c_439_n 0.00377406f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_128 B1 N_A_54_74#_c_439_n 0.0107224f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B1_c_126_n N_A_54_74#_c_429_n 0.00985605f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_130 N_B1_c_126_n N_VGND_c_454_n 6.14068e-19 $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_131 N_B1_c_126_n N_VGND_c_459_n 0.00434272f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_132 N_B1_c_126_n N_VGND_c_463_n 0.00822352f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_133 N_C1_M1006_g N_D1_M1011_g 0.034788f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_134 N_C1_c_158_n N_D1_c_197_n 0.0212265f $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_135 C1 N_D1_c_197_n 5.0774e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_136 N_C1_c_158_n N_D1_c_195_n 0.021434f $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_137 C1 N_D1_c_195_n 0.0128957f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_138 N_C1_c_158_n N_D1_c_196_n 2.00281e-19 $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_139 C1 N_D1_c_196_n 0.0341872f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_140 N_C1_c_158_n N_A_236_368#_c_242_n 5.62853e-19 $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_C1_c_158_n N_A_236_368#_c_243_n 8.2749e-19 $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_C1_c_158_n N_A_236_368#_c_253_n 0.0130996f $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_143 C1 N_A_236_368#_c_253_n 0.0145164f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_144 N_C1_c_158_n N_A_236_368#_c_244_n 0.0111566f $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_145 C1 N_A_236_368#_c_261_n 0.00261116f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_146 N_C1_M1006_g N_A_236_368#_c_234_n 0.00300965f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_147 N_C1_M1006_g N_A_236_368#_c_236_n 7.70038e-19 $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_148 N_C1_c_158_n N_A_236_368#_c_264_n 8.14843e-19 $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_149 C1 N_A_236_368#_c_264_n 0.0254781f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_150 N_C1_c_158_n N_VPWR_c_340_n 0.00833751f $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_151 N_C1_c_158_n N_VPWR_c_341_n 5.65028e-19 $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_152 N_C1_c_158_n N_VPWR_c_348_n 0.00481822f $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_153 N_C1_c_158_n N_VPWR_c_338_n 0.00508379f $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_154 N_C1_M1006_g N_A_54_74#_c_439_n 8.11227e-19 $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_155 N_C1_M1006_g N_A_54_74#_c_429_n 0.00235594f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_156 N_C1_M1006_g N_VGND_c_459_n 0.00461464f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_157 N_C1_M1006_g N_VGND_c_463_n 0.00910941f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_158 N_D1_c_197_n N_A_236_368#_c_244_n 0.00417589f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_D1_c_197_n N_A_236_368#_c_261_n 0.0211153f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_D1_c_195_n N_A_236_368#_c_261_n 0.00174761f $X=2.815 $Y=1.557 $X2=0
+ $Y2=0
cc_161 N_D1_c_196_n N_A_236_368#_c_261_n 0.0254813f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_162 N_D1_M1011_g N_A_236_368#_c_234_n 0.015254f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_163 N_D1_c_195_n N_A_236_368#_c_235_n 5.19479e-19 $X=2.815 $Y=1.557 $X2=0
+ $Y2=0
cc_164 N_D1_c_196_n N_A_236_368#_c_235_n 0.00566599f $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_165 N_D1_M1011_g N_A_236_368#_c_236_n 0.006714f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_166 N_D1_c_195_n N_A_236_368#_c_236_n 0.00435231f $X=2.815 $Y=1.557 $X2=0
+ $Y2=0
cc_167 N_D1_c_196_n N_A_236_368#_c_236_n 0.021921f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_168 N_D1_M1011_g N_A_236_368#_c_237_n 0.00277277f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_169 N_D1_c_195_n N_A_236_368#_c_237_n 0.00116423f $X=2.815 $Y=1.557 $X2=0
+ $Y2=0
cc_170 N_D1_c_196_n N_A_236_368#_c_237_n 0.0150172f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_171 N_D1_c_197_n N_A_236_368#_c_238_n 0.00364448f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_D1_c_195_n N_A_236_368#_c_238_n 4.17225e-19 $X=2.815 $Y=1.557 $X2=0
+ $Y2=0
cc_173 N_D1_c_196_n N_A_236_368#_c_238_n 0.00860662f $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_174 N_D1_M1011_g N_A_236_368#_c_239_n 6.46057e-19 $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_175 N_D1_c_195_n N_A_236_368#_c_239_n 0.0150862f $X=2.815 $Y=1.557 $X2=0
+ $Y2=0
cc_176 N_D1_c_196_n N_A_236_368#_c_239_n 3.56038e-19 $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_177 N_D1_c_197_n N_VPWR_c_341_n 0.0110487f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_178 N_D1_c_197_n N_VPWR_c_348_n 0.00443511f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_179 N_D1_c_197_n N_VPWR_c_338_n 0.00460931f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_180 N_D1_M1011_g N_VGND_c_455_n 0.00373386f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_181 N_D1_M1011_g N_VGND_c_459_n 0.00434272f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_182 N_D1_M1011_g N_VGND_c_463_n 0.00827521f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A_236_368#_c_253_n N_VPWR_M1009_d 0.0179556f $X=2.375 $Y=2.035 $X2=0
+ $Y2=0
cc_184 N_A_236_368#_c_261_n N_VPWR_M1008_d 0.0257579f $X=3.515 $Y=2.035 $X2=0
+ $Y2=0
cc_185 N_A_236_368#_c_238_n N_VPWR_M1008_d 0.00275142f $X=3.6 $Y=1.95 $X2=0
+ $Y2=0
cc_186 N_A_236_368#_c_242_n N_VPWR_c_339_n 0.00823354f $X=1.45 $Y=2.12 $X2=0
+ $Y2=0
cc_187 N_A_236_368#_c_243_n N_VPWR_c_339_n 0.0195335f $X=1.45 $Y=2.695 $X2=0
+ $Y2=0
cc_188 N_A_236_368#_c_243_n N_VPWR_c_340_n 0.0221782f $X=1.45 $Y=2.695 $X2=0
+ $Y2=0
cc_189 N_A_236_368#_c_253_n N_VPWR_c_340_n 0.0249771f $X=2.375 $Y=2.035 $X2=0
+ $Y2=0
cc_190 N_A_236_368#_c_244_n N_VPWR_c_340_n 0.0331292f $X=2.54 $Y=2.375 $X2=0
+ $Y2=0
cc_191 N_A_236_368#_c_240_n N_VPWR_c_341_n 0.017118f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_236_368#_c_244_n N_VPWR_c_341_n 0.0263584f $X=2.54 $Y=2.375 $X2=0
+ $Y2=0
cc_193 N_A_236_368#_c_261_n N_VPWR_c_341_n 0.0604984f $X=3.515 $Y=2.035 $X2=0
+ $Y2=0
cc_194 N_A_236_368#_c_239_n N_VPWR_c_341_n 4.80755e-19 $X=4.245 $Y=1.532 $X2=0
+ $Y2=0
cc_195 N_A_236_368#_c_241_n N_VPWR_c_343_n 0.0261486f $X=4.245 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_236_368#_c_239_n N_VPWR_c_343_n 3.5215e-19 $X=4.245 $Y=1.532 $X2=0
+ $Y2=0
cc_197 N_A_236_368#_c_243_n N_VPWR_c_346_n 0.0097982f $X=1.45 $Y=2.695 $X2=0
+ $Y2=0
cc_198 N_A_236_368#_c_244_n N_VPWR_c_348_n 0.0103753f $X=2.54 $Y=2.375 $X2=0
+ $Y2=0
cc_199 N_A_236_368#_c_240_n N_VPWR_c_349_n 0.00445602f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_236_368#_c_241_n N_VPWR_c_349_n 0.00445602f $X=4.245 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A_236_368#_c_240_n N_VPWR_c_338_n 0.00861719f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_236_368#_c_241_n N_VPWR_c_338_n 0.00860566f $X=4.245 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_236_368#_c_243_n N_VPWR_c_338_n 0.0111907f $X=1.45 $Y=2.695 $X2=0
+ $Y2=0
cc_204 N_A_236_368#_c_244_n N_VPWR_c_338_n 0.0113454f $X=2.54 $Y=2.375 $X2=0
+ $Y2=0
cc_205 N_A_236_368#_c_240_n N_X_c_399_n 0.00261226f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_236_368#_c_241_n N_X_c_399_n 0.00188635f $X=4.245 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_236_368#_c_238_n N_X_c_399_n 0.00559275f $X=3.6 $Y=1.95 $X2=0 $Y2=0
cc_208 N_A_236_368#_c_239_n N_X_c_399_n 0.00697862f $X=4.245 $Y=1.532 $X2=0
+ $Y2=0
cc_209 N_A_236_368#_c_240_n N_X_c_400_n 0.0164541f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_236_368#_c_241_n N_X_c_400_n 0.0109216f $X=4.245 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A_236_368#_M1002_g N_X_c_396_n 0.00104557f $X=3.86 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_236_368#_c_241_n N_X_c_396_n 0.00289345f $X=4.245 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A_236_368#_M1012_g N_X_c_396_n 0.00455396f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_236_368#_c_237_n N_X_c_396_n 0.0293979f $X=3.6 $Y=1.63 $X2=0 $Y2=0
cc_215 N_A_236_368#_c_238_n N_X_c_396_n 0.00661606f $X=3.6 $Y=1.95 $X2=0 $Y2=0
cc_216 N_A_236_368#_c_239_n N_X_c_396_n 0.036292f $X=4.245 $Y=1.532 $X2=0 $Y2=0
cc_217 N_A_236_368#_M1002_g X 0.0122719f $X=3.86 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A_236_368#_M1012_g X 0.00788704f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_236_368#_M1002_g X 0.00479767f $X=3.86 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_236_368#_M1012_g X 0.00327512f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_236_368#_c_237_n X 0.00802092f $X=3.6 $Y=1.63 $X2=0 $Y2=0
cc_222 N_A_236_368#_c_235_n N_VGND_M1002_d 0.00138568f $X=3.515 $Y=1.095 $X2=0
+ $Y2=0
cc_223 N_A_236_368#_c_237_n N_VGND_M1002_d 0.00384491f $X=3.6 $Y=1.63 $X2=0
+ $Y2=0
cc_224 N_A_236_368#_M1002_g N_VGND_c_455_n 0.00634966f $X=3.86 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_236_368#_c_234_n N_VGND_c_455_n 0.032024f $X=3.015 $Y=0.515 $X2=0
+ $Y2=0
cc_226 N_A_236_368#_c_235_n N_VGND_c_455_n 0.00796924f $X=3.515 $Y=1.095 $X2=0
+ $Y2=0
cc_227 N_A_236_368#_c_237_n N_VGND_c_455_n 0.0161682f $X=3.6 $Y=1.63 $X2=0 $Y2=0
cc_228 N_A_236_368#_c_239_n N_VGND_c_455_n 0.00103898f $X=4.245 $Y=1.532 $X2=0
+ $Y2=0
cc_229 N_A_236_368#_M1012_g N_VGND_c_457_n 0.00650681f $X=4.29 $Y=0.74 $X2=0
+ $Y2=0
cc_230 N_A_236_368#_c_234_n N_VGND_c_459_n 0.0145639f $X=3.015 $Y=0.515 $X2=0
+ $Y2=0
cc_231 N_A_236_368#_M1002_g N_VGND_c_460_n 0.00434272f $X=3.86 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_236_368#_M1012_g N_VGND_c_460_n 0.00434272f $X=4.29 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_236_368#_M1002_g N_VGND_c_463_n 0.00825059f $X=3.86 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_236_368#_M1012_g N_VGND_c_463_n 0.00823992f $X=4.29 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_236_368#_c_234_n N_VGND_c_463_n 0.0119984f $X=3.015 $Y=0.515 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_343_n N_X_c_399_n 0.0450694f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_237 N_VPWR_c_341_n N_X_c_400_n 0.0267725f $X=3.52 $Y=2.375 $X2=0 $Y2=0
cc_238 N_VPWR_c_349_n N_X_c_400_n 0.014552f $X=4.355 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_338_n N_X_c_400_n 0.0119791f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_240 X N_VGND_c_455_n 0.0186136f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_241 X N_VGND_c_457_n 0.0293892f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_242 X N_VGND_c_460_n 0.0144922f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_243 X N_VGND_c_463_n 0.0118826f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_244 N_A_54_74#_c_433_n N_VGND_M1010_d 0.0117062f $X=1.39 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_245 N_A_54_74#_c_428_n N_VGND_c_454_n 0.013465f $X=0.485 $Y=0.515 $X2=0 $Y2=0
cc_246 N_A_54_74#_c_433_n N_VGND_c_454_n 0.0279268f $X=1.39 $Y=0.925 $X2=0 $Y2=0
cc_247 N_A_54_74#_c_429_n N_VGND_c_454_n 0.013465f $X=1.555 $Y=0.515 $X2=0 $Y2=0
cc_248 N_A_54_74#_c_428_n N_VGND_c_458_n 0.0146038f $X=0.485 $Y=0.515 $X2=0
+ $Y2=0
cc_249 N_A_54_74#_c_429_n N_VGND_c_459_n 0.0145323f $X=1.555 $Y=0.515 $X2=0
+ $Y2=0
cc_250 N_A_54_74#_c_428_n N_VGND_c_463_n 0.0121018f $X=0.485 $Y=0.515 $X2=0
+ $Y2=0
cc_251 N_A_54_74#_c_433_n N_VGND_c_463_n 0.0114395f $X=1.39 $Y=0.925 $X2=0 $Y2=0
cc_252 N_A_54_74#_c_429_n N_VGND_c_463_n 0.0119861f $X=1.555 $Y=0.515 $X2=0
+ $Y2=0
