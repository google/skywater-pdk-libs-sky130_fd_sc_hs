* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_142_368# B1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.024e+11p pd=2.78e+06u as=7.952e+11p ps=5.9e+06u
M1001 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=6.808e+11p ps=6.28e+06u
M1002 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.255e+11p ps=2.63e+06u
M1003 Y B2 a_142_368# VPB pshort w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=0p ps=0u
M1004 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A1 a_340_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1006 a_340_368# A2 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
