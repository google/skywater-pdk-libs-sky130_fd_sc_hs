* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a222o_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
M1000 VGND C2 a_119_74# VNB nlowvt w=640000u l=150000u
+  ad=9.082e+11p pd=5.52e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_27_390# B1 a_337_390# VPB pshort w=1e+06u l=150000u
+  ad=9.4e+11p pd=7.88e+06u as=7.4e+11p ps=5.48e+06u
M1002 a_337_390# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=8.154e+11p ps=5.8e+06u
M1003 X a_32_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 VPWR A2 a_337_390# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_32_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1006 VGND A2 a_651_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1007 a_651_74# A1 a_32_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=6.848e+11p ps=4.7e+06u
M1008 a_119_74# C1 a_32_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_386_74# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1010 a_32_74# B1 a_386_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_32_74# C1 a_27_390# VPB pshort w=1e+06u l=150000u
+  ad=4.55e+11p pd=2.91e+06u as=0p ps=0u
M1012 a_27_390# C2 a_32_74# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_337_390# B2 a_27_390# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
