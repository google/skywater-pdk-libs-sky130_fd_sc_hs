* File: sky130_fd_sc_hs__o41ai_1.pxi.spice
* Created: Thu Aug 27 21:04:31 2020
* 
x_PM_SKY130_FD_SC_HS__O41AI_1%B1 N_B1_M1009_g N_B1_c_60_n N_B1_M1003_g
+ N_B1_c_57_n N_B1_c_58_n B1 PM_SKY130_FD_SC_HS__O41AI_1%B1
x_PM_SKY130_FD_SC_HS__O41AI_1%A4 N_A4_c_91_n N_A4_M1002_g N_A4_M1008_g A4
+ N_A4_c_93_n PM_SKY130_FD_SC_HS__O41AI_1%A4
x_PM_SKY130_FD_SC_HS__O41AI_1%A3 N_A3_c_131_n N_A3_M1004_g N_A3_M1001_g A3 A3 A3
+ A3 N_A3_c_133_n PM_SKY130_FD_SC_HS__O41AI_1%A3
x_PM_SKY130_FD_SC_HS__O41AI_1%A2 N_A2_M1007_g N_A2_c_173_n N_A2_M1006_g
+ N_A2_c_174_n A2 A2 A2 N_A2_c_177_n A2 PM_SKY130_FD_SC_HS__O41AI_1%A2
x_PM_SKY130_FD_SC_HS__O41AI_1%A1 N_A1_M1000_g N_A1_c_211_n N_A1_M1005_g A1
+ N_A1_c_212_n PM_SKY130_FD_SC_HS__O41AI_1%A1
x_PM_SKY130_FD_SC_HS__O41AI_1%VPWR N_VPWR_M1003_s N_VPWR_M1005_d N_VPWR_c_235_n
+ N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n N_VPWR_c_239_n VPWR
+ N_VPWR_c_240_n N_VPWR_c_234_n PM_SKY130_FD_SC_HS__O41AI_1%VPWR
x_PM_SKY130_FD_SC_HS__O41AI_1%Y N_Y_M1009_s N_Y_M1003_d N_Y_c_268_n N_Y_c_272_n
+ N_Y_c_269_n N_Y_c_280_n N_Y_c_270_n Y N_Y_c_271_n
+ PM_SKY130_FD_SC_HS__O41AI_1%Y
x_PM_SKY130_FD_SC_HS__O41AI_1%A_157_74# N_A_157_74#_M1009_d N_A_157_74#_M1001_d
+ N_A_157_74#_M1000_d N_A_157_74#_c_310_n N_A_157_74#_c_311_n
+ N_A_157_74#_c_312_n N_A_157_74#_c_313_n N_A_157_74#_c_314_n
+ N_A_157_74#_c_315_n N_A_157_74#_c_316_n PM_SKY130_FD_SC_HS__O41AI_1%A_157_74#
x_PM_SKY130_FD_SC_HS__O41AI_1%VGND N_VGND_M1008_d N_VGND_M1007_d N_VGND_c_363_n
+ N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n
+ VGND N_VGND_c_369_n N_VGND_c_370_n PM_SKY130_FD_SC_HS__O41AI_1%VGND
cc_1 VNB N_B1_c_57_n 0.0898718f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_2 VNB N_B1_c_58_n 0.0231039f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.22
cc_3 VNB B1 0.00924172f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A4_c_91_n 0.0269264f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.22
cc_5 VNB N_A4_M1008_g 0.0272905f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.4
cc_6 VNB N_A4_c_93_n 0.00165618f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_7 VNB N_A3_c_131_n 0.0226337f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.22
cc_8 VNB N_A3_M1001_g 0.0259452f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.4
cc_9 VNB N_A3_c_133_n 0.00442043f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_10 VNB N_A2_M1007_g 0.0257812f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.74
cc_11 VNB N_A2_c_173_n 0.0224137f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.4
cc_12 VNB N_A2_c_174_n 0.00484184f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_13 VNB N_A1_M1000_g 0.0348798f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.74
cc_14 VNB N_A1_c_211_n 0.0331637f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.4
cc_15 VNB N_A1_c_212_n 0.015292f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_16 VNB N_VPWR_c_234_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_268_n 0.00273786f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_18 VNB N_Y_c_269_n 0.0036177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_270_n 0.0010381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_271_n 0.0380313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_157_74#_c_310_n 0.00207713f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_22 VNB N_A_157_74#_c_311_n 0.00809218f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_23 VNB N_A_157_74#_c_312_n 0.00541064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_157_74#_c_313_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_157_74#_c_314_n 0.0188655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_157_74#_c_315_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_157_74#_c_316_n 0.00781721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_363_n 0.00977876f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.22
cc_29 VNB N_VGND_c_364_n 0.00970653f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_30 VNB N_VGND_c_365_n 0.0388991f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_31 VNB N_VGND_c_366_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_367_n 0.0191721f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_33 VNB N_VGND_c_368_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_369_n 0.0199471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_370_n 0.215861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B1_c_60_n 0.0188524f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.765
cc_37 VPB N_B1_c_57_n 0.00980037f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.385
cc_38 VPB N_A4_c_91_n 0.027364f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.22
cc_39 VPB N_A4_c_93_n 0.00538051f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_40 VPB N_A3_c_131_n 0.0317629f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.22
cc_41 VPB A3 0.00209573f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.385
cc_42 VPB N_A3_c_133_n 4.05978e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_43 VPB N_A2_c_173_n 0.0327036f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.4
cc_44 VPB N_A2_c_174_n 4.54806e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_45 VPB N_A2_c_177_n 0.00151013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A1_c_211_n 0.0338429f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.4
cc_47 VPB N_A1_c_212_n 0.00936814f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_48 VPB N_VPWR_c_235_n 0.0366602f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.22
cc_49 VPB N_VPWR_c_236_n 0.0303378f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_50 VPB N_VPWR_c_237_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_51 VPB N_VPWR_c_238_n 0.0499688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_239_n 0.0111029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_240_n 0.0682074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_234_n 0.0911385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_Y_c_272_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_56 VPB N_Y_c_270_n 0.00136663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 N_B1_c_60_n N_A4_c_91_n 0.0232424f $X=0.725 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_58 N_B1_c_57_n N_A4_c_91_n 0.02066f $X=0.635 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_59 N_B1_c_57_n N_A4_M1008_g 0.00510291f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_60 N_B1_c_58_n N_A4_M1008_g 0.015975f $X=0.725 $Y=1.22 $X2=0 $Y2=0
cc_61 N_B1_c_57_n N_A4_c_93_n 6.22281e-19 $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_62 N_B1_c_60_n N_VPWR_c_235_n 0.00484854f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_63 N_B1_c_57_n N_VPWR_c_235_n 0.00677105f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_64 B1 N_VPWR_c_235_n 0.0192059f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_B1_c_60_n N_VPWR_c_236_n 0.00592042f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_66 N_B1_c_60_n N_VPWR_c_239_n 0.003296f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_67 N_B1_c_60_n N_VPWR_c_240_n 0.00413917f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_68 N_B1_c_60_n N_VPWR_c_234_n 0.00818241f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_69 N_B1_c_57_n N_Y_c_268_n 0.00705025f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_70 N_B1_c_58_n N_Y_c_268_n 0.00627667f $X=0.725 $Y=1.22 $X2=0 $Y2=0
cc_71 B1 N_Y_c_268_n 0.0124545f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_B1_c_60_n N_Y_c_272_n 0.00464047f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_73 N_B1_c_57_n N_Y_c_269_n 0.0133759f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_74 B1 N_Y_c_269_n 0.0125167f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_B1_c_60_n N_Y_c_280_n 0.00917296f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_76 N_B1_c_60_n N_Y_c_270_n 0.00565543f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_77 N_B1_c_57_n N_Y_c_270_n 0.0127958f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_78 B1 N_Y_c_270_n 0.00143785f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B1_c_57_n N_Y_c_271_n 0.00875781f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_80 N_B1_c_58_n N_Y_c_271_n 0.013685f $X=0.725 $Y=1.22 $X2=0 $Y2=0
cc_81 B1 N_Y_c_271_n 0.0273814f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_B1_c_58_n N_A_157_74#_c_310_n 0.00464354f $X=0.725 $Y=1.22 $X2=0 $Y2=0
cc_83 N_B1_c_58_n N_A_157_74#_c_312_n 0.00131473f $X=0.725 $Y=1.22 $X2=0 $Y2=0
cc_84 N_B1_c_58_n N_VGND_c_365_n 0.00303976f $X=0.725 $Y=1.22 $X2=0 $Y2=0
cc_85 N_B1_c_58_n N_VGND_c_370_n 0.00404638f $X=0.725 $Y=1.22 $X2=0 $Y2=0
cc_86 N_A4_c_91_n N_A3_c_131_n 0.0646419f $X=1.225 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_87 N_A4_c_93_n N_A3_c_131_n 6.85744e-19 $X=1.22 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_88 N_A4_M1008_g N_A3_M1001_g 0.0248295f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A4_c_91_n A3 0.0107861f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A4_c_93_n A3 0.0077832f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A4_c_91_n N_A3_c_133_n 0.00201946f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A4_c_93_n N_A3_c_133_n 0.0253181f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_93 N_A4_c_91_n N_VPWR_c_236_n 5.20254e-19 $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A4_c_91_n N_VPWR_c_240_n 0.00445602f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A4_c_91_n N_VPWR_c_234_n 0.00859297f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A4_M1008_g N_Y_c_268_n 9.38286e-19 $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A4_c_91_n N_Y_c_272_n 0.0132887f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A4_c_91_n N_Y_c_269_n 9.98351e-19 $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A4_c_93_n N_Y_c_269_n 0.0131895f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A4_c_91_n N_Y_c_280_n 0.00305835f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A4_c_93_n N_Y_c_280_n 0.00688138f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A4_c_91_n N_Y_c_270_n 0.00429768f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A4_c_93_n N_Y_c_270_n 0.0199517f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A4_M1008_g N_Y_c_271_n 3.37387e-19 $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A4_M1008_g N_A_157_74#_c_310_n 0.00959047f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A4_c_91_n N_A_157_74#_c_311_n 3.80672e-19 $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A4_M1008_g N_A_157_74#_c_311_n 0.0118537f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A4_c_93_n N_A_157_74#_c_311_n 0.0132954f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A4_c_91_n N_A_157_74#_c_312_n 9.78174e-19 $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A4_M1008_g N_A_157_74#_c_312_n 0.00154351f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A4_c_93_n N_A_157_74#_c_312_n 0.0127466f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_112 N_A4_M1008_g N_A_157_74#_c_313_n 8.69432e-19 $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A4_M1008_g N_VGND_c_363_n 0.00633237f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A4_M1008_g N_VGND_c_365_n 0.00434272f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A4_M1008_g N_VGND_c_370_n 0.00822486f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A3_M1001_g N_A2_M1007_g 0.0199862f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A3_c_131_n N_A2_c_173_n 0.0563226f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_118 A3 N_A2_c_173_n 0.00101838f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_119 N_A3_c_133_n N_A2_c_173_n 3.62017e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A3_c_131_n N_A2_c_174_n 0.00114507f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A3_c_133_n N_A2_c_174_n 0.0269386f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A3_c_131_n A2 0.00378834f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A3_c_131_n N_A2_c_177_n 0.00112827f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_124 A3 N_A2_c_177_n 0.00918143f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A3_c_131_n N_VPWR_c_240_n 0.00303293f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_126 A3 N_VPWR_c_240_n 0.0060786f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A3_c_131_n N_VPWR_c_234_n 0.00373561f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_128 A3 N_VPWR_c_234_n 0.00720215f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A3_c_131_n N_Y_c_272_n 4.19885e-19 $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A3_c_131_n N_Y_c_280_n 9.08111e-19 $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_131 A3 N_Y_c_280_n 0.0368511f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_132 A3 A_260_368# 0.0134616f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_133 N_A3_M1001_g N_A_157_74#_c_310_n 8.64759e-19 $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A3_c_131_n N_A_157_74#_c_311_n 0.00364765f $X=1.715 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A3_M1001_g N_A_157_74#_c_311_n 0.0118588f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A3_c_133_n N_A_157_74#_c_311_n 0.0241717f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A3_M1001_g N_A_157_74#_c_313_n 0.00988375f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A3_c_131_n N_A_157_74#_c_316_n 9.31826e-19 $X=1.715 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A3_M1001_g N_A_157_74#_c_316_n 0.00155819f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A3_c_133_n N_A_157_74#_c_316_n 0.00536895f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A3_M1001_g N_VGND_c_363_n 0.00781129f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A3_M1001_g N_VGND_c_367_n 0.00434272f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A3_M1001_g N_VGND_c_370_n 0.00821853f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A2_M1007_g N_A1_M1000_g 0.0260254f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A2_c_173_n N_A1_c_211_n 0.0553536f $X=2.285 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A2_c_174_n N_A1_c_211_n 0.00127309f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A2_c_177_n N_A1_c_211_n 0.00595528f $X=2.17 $Y=1.92 $X2=0 $Y2=0
cc_148 N_A2_c_173_n N_A1_c_212_n 7.4401e-19 $X=2.285 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A2_c_174_n N_A1_c_212_n 0.0169052f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A2_c_177_n N_A1_c_212_n 0.0029171f $X=2.17 $Y=1.92 $X2=0 $Y2=0
cc_151 N_A2_c_173_n N_VPWR_c_240_n 0.00372889f $X=2.285 $Y=1.765 $X2=0 $Y2=0
cc_152 A2 N_VPWR_c_240_n 0.00687333f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_153 N_A2_c_173_n N_VPWR_c_234_n 0.00610745f $X=2.285 $Y=1.765 $X2=0 $Y2=0
cc_154 A2 N_VPWR_c_234_n 0.00822835f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_155 A2 A_358_368# 0.0149411f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_156 N_A2_c_177_n A_358_368# 9.30302e-19 $X=2.17 $Y=1.92 $X2=-0.19 $Y2=-0.245
cc_157 N_A2_M1007_g N_A_157_74#_c_313_n 0.00966073f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1007_g N_A_157_74#_c_314_n 0.0117984f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_c_173_n N_A_157_74#_c_314_n 0.00411108f $X=2.285 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A2_c_174_n N_A_157_74#_c_314_n 0.0224209f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A2_M1007_g N_A_157_74#_c_315_n 6.28869e-19 $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A2_M1007_g N_A_157_74#_c_316_n 0.00155819f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A2_c_174_n N_A_157_74#_c_316_n 0.00818793f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A2_M1007_g N_VGND_c_364_n 0.00622602f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A2_M1007_g N_VGND_c_367_n 0.00434272f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A2_M1007_g N_VGND_c_370_n 0.0082141f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_c_211_n N_VPWR_c_238_n 0.0275375f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A1_c_212_n N_VPWR_c_238_n 0.0211526f $X=2.975 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A1_c_211_n N_VPWR_c_240_n 0.00461464f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A1_c_211_n N_VPWR_c_234_n 0.009135f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A1_M1000_g N_A_157_74#_c_313_n 6.28869e-19 $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A1_M1000_g N_A_157_74#_c_314_n 0.0153182f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A1_c_211_n N_A_157_74#_c_314_n 0.00177898f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A1_c_212_n N_A_157_74#_c_314_n 0.0344691f $X=2.975 $Y=1.515 $X2=0 $Y2=0
cc_175 N_A1_M1000_g N_A_157_74#_c_315_n 0.0103339f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_M1000_g N_VGND_c_364_n 0.00622602f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A1_M1000_g N_VGND_c_369_n 0.00434272f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A1_M1000_g N_VGND_c_370_n 0.00825053f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_179 N_VPWR_c_239_n N_Y_c_272_n 0.0141382f $X=0.495 $Y=2.815 $X2=0 $Y2=0
cc_180 N_VPWR_c_240_n N_Y_c_272_n 0.0145938f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VPWR_c_234_n N_Y_c_272_n 0.0120466f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_182 N_VPWR_c_235_n N_Y_c_270_n 0.0236075f $X=0.455 $Y=1.985 $X2=0 $Y2=0
cc_183 N_Y_c_271_n N_A_157_74#_c_310_n 0.0505664f $X=0.495 $Y=0.515 $X2=0 $Y2=0
cc_184 N_Y_c_268_n N_A_157_74#_c_312_n 0.0129299f $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_185 N_Y_c_271_n N_VGND_c_365_n 0.0284523f $X=0.495 $Y=0.515 $X2=0 $Y2=0
cc_186 N_Y_c_271_n N_VGND_c_370_n 0.0232443f $X=0.495 $Y=0.515 $X2=0 $Y2=0
cc_187 N_A_157_74#_c_311_n N_VGND_M1008_d 0.00378075f $X=1.89 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_157_74#_c_314_n N_VGND_M1007_d 0.00358162f $X=2.89 $Y=1.095 $X2=0
+ $Y2=0
cc_189 N_A_157_74#_c_310_n N_VGND_c_363_n 0.0184106f $X=1.04 $Y=0.515 $X2=0
+ $Y2=0
cc_190 N_A_157_74#_c_311_n N_VGND_c_363_n 0.0257907f $X=1.89 $Y=1.095 $X2=0
+ $Y2=0
cc_191 N_A_157_74#_c_313_n N_VGND_c_363_n 0.0356652f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_192 N_A_157_74#_c_313_n N_VGND_c_364_n 0.0191765f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_193 N_A_157_74#_c_314_n N_VGND_c_364_n 0.0248957f $X=2.89 $Y=1.095 $X2=0
+ $Y2=0
cc_194 N_A_157_74#_c_315_n N_VGND_c_364_n 0.0191765f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
cc_195 N_A_157_74#_c_310_n N_VGND_c_365_n 0.0109942f $X=1.04 $Y=0.515 $X2=0
+ $Y2=0
cc_196 N_A_157_74#_c_313_n N_VGND_c_367_n 0.0144922f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_197 N_A_157_74#_c_315_n N_VGND_c_369_n 0.0145639f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
cc_198 N_A_157_74#_c_310_n N_VGND_c_370_n 0.00904371f $X=1.04 $Y=0.515 $X2=0
+ $Y2=0
cc_199 N_A_157_74#_c_313_n N_VGND_c_370_n 0.0118826f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_200 N_A_157_74#_c_315_n N_VGND_c_370_n 0.0119984f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
