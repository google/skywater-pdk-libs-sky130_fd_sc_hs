* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
M1000 Y A1 a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=1.0767e+12p pd=1.031e+07u as=8.917e+11p ps=8.33e+06u
M1001 a_114_85# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_478_368# S VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=1.4448e+12p pd=1.154e+07u as=2.5466e+12p ps=1.762e+07u
M1003 a_478_368# A0 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.792e+12p ps=1.44e+07u
M1004 a_478_368# S VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_475_85# A0 Y VNB nlowvt w=740000u l=150000u
+  ad=8.806e+11p pd=8.3e+06u as=0p ps=0u
M1006 VPWR a_1030_268# a_116_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.4336e+12p ps=1.152e+07u
M1007 VPWR S a_478_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_114_85# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.795e+12p ps=1.331e+07u
M1009 VPWR S a_478_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1030_268# S VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1011 a_475_85# a_1030_268# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_1030_268# a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_114_85# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR S a_1030_268# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_116_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_116_368# A1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_114_85# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_116_368# A1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A1 a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1030_268# S VGND VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1021 a_116_368# a_1030_268# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A1 a_116_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_478_368# A0 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y A0 a_478_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1030_268# a_116_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND S a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A0 a_478_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_1030_268# a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_116_368# a_1030_268# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND S a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_475_85# a_1030_268# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y A0 a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y A0 a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_475_85# A0 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
