* File: sky130_fd_sc_hs__sdfrtn_1.spice
* Created: Tue Sep  1 20:22:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfrtn_1.pex.spice"
.subckt sky130_fd_sc_hs__sdfrtn_1  VNB VPB SCE D SCD RESET_B CLK_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK_N	CLK_N
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1037 N_VGND_M1037_d N_SCE_M1037_g N_A_27_88#_M1037_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1491 AS=0.1197 PD=1.55 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 noxref_25 N_A_27_88#_M1013_g N_noxref_24_M1013_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1014 N_A_284_464#_M1014_d N_D_M1014_g noxref_25 VNB NLOWVT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=0.98 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1003 noxref_26 N_SCE_M1003_g N_A_284_464#_M1014_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1176 PD=0.66 PS=0.98 NRD=18.564 NRS=39.996 M=1 R=2.8 SA=75001.3
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1033 N_noxref_24_M1033_d N_SCD_M1033_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.0609 AS=0.0504 PD=0.71 PS=0.66 NRD=1.428 NRS=18.564 M=1 R=2.8 SA=75001.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_RESET_B_M1022_g N_noxref_24_M1033_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.161981 AS=0.0609 PD=1.14052 PS=0.71 NRD=94.476 NRS=1.428 M=1 R=2.8
+ SA=75002.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1009 N_A_854_74#_M1009_d N_CLK_N_M1009_g N_VGND_M1022_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.285394 PD=2.05 PS=2.00948 NRD=0 NRS=53.616 M=1 R=4.93333
+ SA=75001.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_1074_88#_M1015_d N_A_854_74#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.3899 PD=2.05 PS=2.88 NRD=0 NRS=76.512 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_A_1272_131#_M1027_d N_A_1074_88#_M1027_g N_A_284_464#_M1027_s VNB
+ NLOWVT L=0.15 W=0.42 AD=0.11445 AS=0.1197 PD=0.965 PS=1.41 NRD=72.852 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1023 A_1411_131# N_A_854_74#_M1023_g N_A_1272_131#_M1027_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.11445 PD=0.66 PS=0.965 NRD=18.564 NRS=2.856 M=1 R=2.8
+ SA=75000.9 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1034 A_1489_131# N_A_1429_308#_M1034_g A_1411_131# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_RESET_B_M1018_g A_1489_131# VNB NLOWVT L=0.15 W=0.42
+ AD=0.129972 AS=0.0504 PD=1.11736 PS=0.66 NRD=72.696 NRS=18.564 M=1 R=2.8
+ SA=75001.7 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1035 N_A_1429_308#_M1035_d N_A_1272_131#_M1035_g N_VGND_M1018_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1792 AS=0.198053 PD=1.2 PS=1.70264 NRD=26.244 NRS=47.7 M=1
+ R=4.26667 SA=75001.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1039 N_A_1827_144#_M1039_d N_A_854_74#_M1039_g N_A_1429_308#_M1035_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.377751 AS=0.1792 PD=2.57208 PS=1.2 NRD=100.356
+ NRS=26.244 M=1 R=4.26667 SA=75002 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1028 A_2073_74# N_A_1074_88#_M1028_g N_A_1827_144#_M1039_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0525 AS=0.247899 PD=0.67 PS=1.68792 NRD=19.992 NRS=24.276 M=1
+ R=2.8 SA=75001.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_2087_410#_M1001_g A_2073_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0861 AS=0.0525 PD=0.83 PS=0.67 NRD=17.136 NRS=19.992 M=1 R=2.8 SA=75001.9
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 A_2265_74# N_RESET_B_M1004_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0861 PD=0.66 PS=0.83 NRD=18.564 NRS=19.992 M=1 R=2.8 SA=75002.4
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_A_2087_410#_M1005_d N_A_1827_144#_M1005_g A_2265_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.21 AS=0.0504 PD=1.84 PS=0.66 NRD=30 NRS=18.564 M=1 R=2.8
+ SA=75002.8 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1827_144#_M1029_g N_A_2492_424#_M1029_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=25.632 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1010 N_Q_M1010_d N_A_2492_424#_M1010_g N_VGND_M1029_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VPWR_M1016_d N_SCE_M1016_g N_A_27_88#_M1016_s VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.1888 PD=0.94 PS=1.87 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75003 A=0.096 P=1.58 MULT=1
MM1017 A_206_464# N_SCE_M1017_g N_VPWR_M1016_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.096 PD=0.88 PS=0.94 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_284_464#_M1002_d N_D_M1002_g A_206_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.2512 AS=0.0768 PD=1.425 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75001.1 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1036 A_471_464# N_A_27_88#_M1036_g N_A_284_464#_M1002_d VPB PSHORT L=0.15
+ W=0.64 AD=0.0768 AS=0.2512 PD=0.88 PS=1.425 NRD=19.9955 NRS=3.0732 M=1
+ R=4.26667 SA=75002 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_SCD_M1006_g A_471_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.184475 AS=0.0768 PD=1.345 PS=0.88 NRD=71.7868 NRS=19.9955 M=1 R=4.26667
+ SA=75002.4 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1012 N_A_284_464#_M1012_d N_RESET_B_M1012_g N_VPWR_M1006_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1888 AS=0.184475 PD=1.87 PS=1.345 NRD=3.0732 NRS=71.7868 M=1
+ R=4.26667 SA=75003 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1038 N_A_854_74#_M1038_d N_CLK_N_M1038_g N_VPWR_M1038_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.4144 PD=2.83 PS=2.98 NRD=1.7533 NRS=14.9326 M=1
+ R=7.46667 SA=75000.3 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1026 N_A_1074_88#_M1026_d N_A_854_74#_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1020 N_A_1272_131#_M1020_d N_A_854_74#_M1020_g N_A_284_464#_M1020_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1024 A_1384_508# N_A_1074_88#_M1024_g N_A_1272_131#_M1020_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.063 PD=0.66 PS=0.72 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_1429_308#_M1007_g A_1384_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.0504 PD=0.72 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_A_1272_131#_M1011_d N_RESET_B_M1011_g N_VPWR_M1007_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1239 AS=0.063 PD=1.43 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_1429_308#_M1025_d N_A_1272_131#_M1025_g N_VPWR_M1025_s VPB PSHORT
+ L=0.15 W=1 AD=0.3925 AS=0.285 PD=1.785 PS=2.57 NRD=11.8003 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1000 N_A_1827_144#_M1000_d N_A_1074_88#_M1000_g N_A_1429_308#_M1025_d VPB
+ PSHORT L=0.15 W=1 AD=0.220282 AS=0.3925 PD=1.92254 PS=1.785 NRD=5.5751
+ NRS=1.9503 M=1 R=6.66667 SA=75001.1 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1031 A_2042_508# N_A_854_74#_M1031_g N_A_1827_144#_M1000_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0546 AS=0.0925183 PD=0.68 PS=0.807465 NRD=35.1645 NRS=23.443 M=1
+ R=2.8 SA=75001.7 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_2087_410#_M1021_g A_2042_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.13125 AS=0.0546 PD=1.045 PS=0.68 NRD=68.0044 NRS=35.1645 M=1 R=2.8
+ SA=75002.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1030 N_A_2087_410#_M1030_d N_RESET_B_M1030_g N_VPWR_M1021_d VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.13125 PD=0.72 PS=1.045 NRD=4.6886 NRS=93.7917 M=1 R=2.8
+ SA=75002.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_1827_144#_M1032_g N_A_2087_410#_M1030_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.1449 AS=0.063 PD=1.53 PS=0.72 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75003.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_1827_144#_M1008_g N_A_2492_424#_M1008_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1956 AS=0.2478 PD=1.32857 PS=2.27 NRD=22.261 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1019 N_Q_M1019_d N_A_2492_424#_M1019_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1.12
+ AD=0.336 AS=0.2608 PD=2.84 PS=1.77143 NRD=2.6201 NRS=9.6727 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=26.1504 P=32.56
*
.include "sky130_fd_sc_hs__sdfrtn_1.pxi.spice"
*
.ends
*
*
