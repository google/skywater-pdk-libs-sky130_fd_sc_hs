* File: sky130_fd_sc_hs__mux4_2.pxi.spice
* Created: Tue Sep  1 20:08:17 2020
* 
x_PM_SKY130_FD_SC_HS__MUX4_2%S0 N_S0_M1001_g N_S0_c_165_n N_S0_c_183_n
+ N_S0_M1007_g N_S0_M1010_g N_S0_c_167_n N_S0_M1020_g N_S0_M1016_g N_S0_c_168_n
+ N_S0_M1022_g N_S0_c_283_p N_S0_c_206_p N_S0_c_319_p N_S0_c_207_p N_S0_c_169_n
+ N_S0_c_170_n N_S0_c_171_n N_S0_c_172_n N_S0_c_173_n N_S0_c_174_n N_S0_c_175_n
+ N_S0_c_176_n N_S0_c_177_n S0 N_S0_c_179_n N_S0_c_180_n N_S0_c_181_n
+ PM_SKY130_FD_SC_HS__MUX4_2%S0
x_PM_SKY130_FD_SC_HS__MUX4_2%A1 N_A1_M1013_g N_A1_c_329_n N_A1_M1002_g A1
+ PM_SKY130_FD_SC_HS__MUX4_2%A1
x_PM_SKY130_FD_SC_HS__MUX4_2%A_31_94# N_A_31_94#_M1001_s N_A_31_94#_M1007_s
+ N_A_31_94#_c_359_n N_A_31_94#_M1000_g N_A_31_94#_M1014_g N_A_31_94#_c_361_n
+ N_A_31_94#_M1015_g N_A_31_94#_M1005_g N_A_31_94#_c_369_n N_A_31_94#_c_363_n
+ N_A_31_94#_c_399_n N_A_31_94#_c_370_n N_A_31_94#_c_402_n N_A_31_94#_c_371_n
+ N_A_31_94#_c_372_n N_A_31_94#_c_373_n N_A_31_94#_c_364_n N_A_31_94#_c_365_n
+ N_A_31_94#_c_366_n PM_SKY130_FD_SC_HS__MUX4_2%A_31_94#
x_PM_SKY130_FD_SC_HS__MUX4_2%A0 N_A0_M1023_g N_A0_c_480_n N_A0_c_481_n
+ N_A0_c_482_n N_A0_M1004_g A0 PM_SKY130_FD_SC_HS__MUX4_2%A0
x_PM_SKY130_FD_SC_HS__MUX4_2%A3 N_A3_M1019_g N_A3_c_519_n N_A3_M1003_g A3
+ PM_SKY130_FD_SC_HS__MUX4_2%A3
x_PM_SKY130_FD_SC_HS__MUX4_2%A2 N_A2_M1011_g N_A2_c_552_n N_A2_c_557_n
+ N_A2_M1026_g A2 A2 N_A2_c_554_n N_A2_c_555_n PM_SKY130_FD_SC_HS__MUX4_2%A2
x_PM_SKY130_FD_SC_HS__MUX4_2%A_1500_94# N_A_1500_94#_M1008_s
+ N_A_1500_94#_M1018_s N_A_1500_94#_c_596_n N_A_1500_94#_M1006_g
+ N_A_1500_94#_c_601_n N_A_1500_94#_M1017_g N_A_1500_94#_c_597_n
+ N_A_1500_94#_c_598_n N_A_1500_94#_c_603_n N_A_1500_94#_c_599_n
+ N_A_1500_94#_c_600_n PM_SKY130_FD_SC_HS__MUX4_2%A_1500_94#
x_PM_SKY130_FD_SC_HS__MUX4_2%S1 N_S1_M1009_g N_S1_c_651_n N_S1_M1012_g
+ N_S1_c_652_n N_S1_c_653_n N_S1_M1008_g N_S1_c_655_n N_S1_c_656_n N_S1_c_660_n
+ N_S1_M1018_g S1 PM_SKY130_FD_SC_HS__MUX4_2%S1
x_PM_SKY130_FD_SC_HS__MUX4_2%A_1429_74# N_A_1429_74#_M1009_d
+ N_A_1429_74#_M1012_d N_A_1429_74#_c_728_n N_A_1429_74#_M1021_g
+ N_A_1429_74#_c_736_n N_A_1429_74#_M1024_g N_A_1429_74#_c_729_n
+ N_A_1429_74#_M1025_g N_A_1429_74#_c_737_n N_A_1429_74#_M1027_g
+ N_A_1429_74#_c_730_n N_A_1429_74#_c_731_n N_A_1429_74#_c_732_n
+ N_A_1429_74#_c_740_n N_A_1429_74#_c_733_n N_A_1429_74#_c_741_n
+ N_A_1429_74#_c_734_n N_A_1429_74#_c_742_n N_A_1429_74#_c_735_n
+ PM_SKY130_FD_SC_HS__MUX4_2%A_1429_74#
x_PM_SKY130_FD_SC_HS__MUX4_2%VPWR N_VPWR_M1007_d N_VPWR_M1004_d N_VPWR_M1026_d
+ N_VPWR_M1018_d N_VPWR_M1027_s N_VPWR_c_833_n N_VPWR_c_834_n N_VPWR_c_835_n
+ N_VPWR_c_836_n N_VPWR_c_837_n N_VPWR_c_838_n N_VPWR_c_839_n N_VPWR_c_840_n
+ N_VPWR_c_841_n N_VPWR_c_842_n N_VPWR_c_843_n VPWR N_VPWR_c_844_n
+ N_VPWR_c_845_n N_VPWR_c_846_n N_VPWR_c_847_n N_VPWR_c_832_n
+ PM_SKY130_FD_SC_HS__MUX4_2%VPWR
x_PM_SKY130_FD_SC_HS__MUX4_2%A_333_74# N_A_333_74#_M1010_d N_A_333_74#_M1006_d
+ N_A_333_74#_M1000_d N_A_333_74#_M1012_s N_A_333_74#_c_946_n
+ N_A_333_74#_c_937_n N_A_333_74#_c_972_n N_A_333_74#_c_975_n
+ N_A_333_74#_c_997_n N_A_333_74#_c_938_n N_A_333_74#_c_939_n
+ N_A_333_74#_c_933_n N_A_333_74#_c_934_n N_A_333_74#_c_935_n
+ N_A_333_74#_c_941_n N_A_333_74#_c_942_n N_A_333_74#_c_936_n
+ N_A_333_74#_c_944_n PM_SKY130_FD_SC_HS__MUX4_2%A_333_74#
x_PM_SKY130_FD_SC_HS__MUX4_2%A_909_74# N_A_909_74#_M1016_d N_A_909_74#_M1009_s
+ N_A_909_74#_M1015_d N_A_909_74#_M1017_d N_A_909_74#_c_1078_n
+ N_A_909_74#_c_1065_n N_A_909_74#_c_1072_n N_A_909_74#_c_1066_n
+ N_A_909_74#_c_1098_n N_A_909_74#_c_1073_n N_A_909_74#_c_1074_n
+ N_A_909_74#_c_1067_n N_A_909_74#_c_1068_n N_A_909_74#_c_1069_n
+ N_A_909_74#_c_1096_n N_A_909_74#_c_1070_n N_A_909_74#_c_1076_n
+ N_A_909_74#_c_1071_n PM_SKY130_FD_SC_HS__MUX4_2%A_909_74#
x_PM_SKY130_FD_SC_HS__MUX4_2%X N_X_M1021_d N_X_M1024_d X X X X X X X X
+ PM_SKY130_FD_SC_HS__MUX4_2%X
x_PM_SKY130_FD_SC_HS__MUX4_2%VGND N_VGND_M1001_d N_VGND_M1023_d N_VGND_M1011_d
+ N_VGND_M1008_d N_VGND_M1025_s N_VGND_c_1222_n N_VGND_c_1223_n N_VGND_c_1224_n
+ N_VGND_c_1225_n N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n
+ N_VGND_c_1229_n N_VGND_c_1230_n N_VGND_c_1231_n VGND N_VGND_c_1232_n
+ N_VGND_c_1233_n N_VGND_c_1234_n N_VGND_c_1235_n N_VGND_c_1236_n
+ N_VGND_c_1237_n PM_SKY130_FD_SC_HS__MUX4_2%VGND
cc_1 VNB N_S0_c_165_n 0.00667767f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.795
cc_2 VNB N_S0_M1010_g 0.0223899f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=0.74
cc_3 VNB N_S0_c_167_n 0.0256351f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=1.885
cc_4 VNB N_S0_c_168_n 0.0259677f $X=-0.19 $Y=-0.245 $X2=5.685 $Y2=1.885
cc_5 VNB N_S0_c_169_n 0.00286293f $X=-0.19 $Y=-0.245 $X2=2.94 $Y2=1.615
cc_6 VNB N_S0_c_170_n 0.0357364f $X=-0.19 $Y=-0.245 $X2=4.395 $Y2=1.195
cc_7 VNB N_S0_c_171_n 0.023949f $X=-0.19 $Y=-0.245 $X2=5.475 $Y2=1.195
cc_8 VNB N_S0_c_172_n 0.00237512f $X=-0.19 $Y=-0.245 $X2=5.64 $Y2=1.585
cc_9 VNB N_S0_c_173_n 0.0317907f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.195
cc_10 VNB N_S0_c_174_n 0.0351747f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.425
cc_11 VNB N_S0_c_175_n 0.0027148f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.195
cc_12 VNB N_S0_c_176_n 0.00555302f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.195
cc_13 VNB N_S0_c_177_n 0.037993f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.385
cc_14 VNB S0 0.0102619f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_15 VNB N_S0_c_179_n 0.0351679f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_16 VNB N_S0_c_180_n 0.022866f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.22
cc_17 VNB N_S0_c_181_n 0.0181052f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.22
cc_18 VNB N_A1_M1013_g 0.0299746f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.79
cc_19 VNB N_A1_c_329_n 0.0174636f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.795
cc_20 VNB A1 0.00539029f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.46
cc_21 VNB N_A_31_94#_c_359_n 0.0313605f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.46
cc_22 VNB N_A_31_94#_M1014_g 0.042397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_31_94#_c_361_n 0.0194956f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=2.46
cc_24 VNB N_A_31_94#_M1005_g 0.0381472f $X=-0.19 $Y=-0.245 $X2=5.685 $Y2=1.885
cc_25 VNB N_A_31_94#_c_363_n 0.0210344f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.28
cc_26 VNB N_A_31_94#_c_364_n 0.00699674f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.195
cc_27 VNB N_A_31_94#_c_365_n 0.00649887f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.385
cc_28 VNB N_A_31_94#_c_366_n 0.0299914f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.55
cc_29 VNB N_A0_M1023_g 0.0242281f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.79
cc_30 VNB N_A0_c_480_n 0.0186106f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.795
cc_31 VNB N_A0_c_481_n 0.0126854f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.885
cc_32 VNB N_A0_c_482_n 0.00249175f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.46
cc_33 VNB A0 0.00301611f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=0.74
cc_34 VNB N_A3_M1019_g 0.0302618f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.79
cc_35 VNB N_A3_c_519_n 0.0180435f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.795
cc_36 VNB A3 0.00614143f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.46
cc_37 VNB N_A2_c_552_n 0.00579376f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.795
cc_38 VNB A2 0.00748937f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.26
cc_39 VNB N_A2_c_554_n 0.0375536f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=2.46
cc_40 VNB N_A2_c_555_n 0.0242171f $X=-0.19 $Y=-0.245 $X2=4.47 $Y2=1.22
cc_41 VNB N_A_1500_94#_c_596_n 0.0205391f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.46
cc_42 VNB N_A_1500_94#_c_597_n 0.0106693f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=2.46
cc_43 VNB N_A_1500_94#_c_598_n 0.0079758f $X=-0.19 $Y=-0.245 $X2=5.685 $Y2=1.885
cc_44 VNB N_A_1500_94#_c_599_n 0.00129826f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=0.59
cc_45 VNB N_A_1500_94#_c_600_n 0.0448895f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.11
cc_46 VNB N_S1_M1009_g 0.0290609f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.55
cc_47 VNB N_S1_c_651_n 0.0239793f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.795
cc_48 VNB N_S1_c_652_n 0.121123f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.46
cc_49 VNB N_S1_c_653_n 0.012589f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.26
cc_50 VNB N_S1_M1008_g 0.0319136f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=1.885
cc_51 VNB N_S1_c_655_n 0.00770192f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=2.46
cc_52 VNB N_S1_c_656_n 0.0129905f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=2.46
cc_53 VNB S1 0.00428476f $X=-0.19 $Y=-0.245 $X2=5.685 $Y2=2.46
cc_54 VNB N_A_1429_74#_c_728_n 0.017253f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.46
cc_55 VNB N_A_1429_74#_c_729_n 0.0188588f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=1.885
cc_56 VNB N_A_1429_74#_c_730_n 0.036345f $X=-0.19 $Y=-0.245 $X2=5.685 $Y2=1.885
cc_57 VNB N_A_1429_74#_c_731_n 0.0502811f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=0.59
cc_58 VNB N_A_1429_74#_c_732_n 0.0224813f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=0.505
cc_59 VNB N_A_1429_74#_c_733_n 0.00594835f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.615
cc_60 VNB N_A_1429_74#_c_734_n 0.00358595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1429_74#_c_735_n 0.00213054f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.425
cc_62 VNB N_VPWR_c_832_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_333_74#_c_933_n 0.00779776f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.28
cc_64 VNB N_A_333_74#_c_934_n 0.00419076f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.615
cc_65 VNB N_A_333_74#_c_935_n 0.00961107f $X=-0.19 $Y=-0.245 $X2=2.94 $Y2=1.615
cc_66 VNB N_A_333_74#_c_936_n 0.00416275f $X=-0.19 $Y=-0.245 $X2=5.61 $Y2=1.585
cc_67 VNB N_A_909_74#_c_1065_n 0.0104114f $X=-0.19 $Y=-0.245 $X2=4.47 $Y2=0.74
cc_68 VNB N_A_909_74#_c_1066_n 0.00708214f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.11
cc_69 VNB N_A_909_74#_c_1067_n 0.00810674f $X=-0.19 $Y=-0.245 $X2=4.395
+ $Y2=1.195
cc_70 VNB N_A_909_74#_c_1068_n 0.00389352f $X=-0.19 $Y=-0.245 $X2=4.725
+ $Y2=1.195
cc_71 VNB N_A_909_74#_c_1069_n 0.00475336f $X=-0.19 $Y=-0.245 $X2=5.61 $Y2=1.585
cc_72 VNB N_A_909_74#_c_1070_n 3.81574e-19 $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.195
cc_73 VNB N_A_909_74#_c_1071_n 0.00515798f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.385
cc_74 VNB X 0.00279061f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.46
cc_75 VNB N_VGND_c_1222_n 0.0103581f $X=-0.19 $Y=-0.245 $X2=4.47 $Y2=0.74
cc_76 VNB N_VGND_c_1223_n 0.00825158f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=0.505
cc_77 VNB N_VGND_c_1224_n 0.00906639f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.28
cc_78 VNB N_VGND_c_1225_n 0.0138034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1226_n 0.0117944f $X=-0.19 $Y=-0.245 $X2=3.105 $Y2=1.195
cc_80 VNB N_VGND_c_1227_n 0.0556926f $X=-0.19 $Y=-0.245 $X2=4.725 $Y2=1.195
cc_81 VNB N_VGND_c_1228_n 0.0260969f $X=-0.19 $Y=-0.245 $X2=5.64 $Y2=1.585
cc_82 VNB N_VGND_c_1229_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=5.64 $Y2=1.585
cc_83 VNB N_VGND_c_1230_n 0.0657879f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.195
cc_84 VNB N_VGND_c_1231_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.195
cc_85 VNB N_VGND_c_1232_n 0.0616371f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.385
cc_86 VNB N_VGND_c_1233_n 0.0685518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1234_n 0.0197463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1235_n 0.00904775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1236_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1237_n 0.586934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VPB N_S0_c_165_n 0.00828485f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.795
cc_92 VPB N_S0_c_183_n 0.0290863f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.885
cc_93 VPB N_S0_c_167_n 0.0377368f $X=-0.19 $Y=1.66 $X2=3.015 $Y2=1.885
cc_94 VPB N_S0_c_168_n 0.0369031f $X=-0.19 $Y=1.66 $X2=5.685 $Y2=1.885
cc_95 VPB N_S0_c_169_n 6.81649e-19 $X=-0.19 $Y=1.66 $X2=2.94 $Y2=1.615
cc_96 VPB N_S0_c_172_n 0.00120129f $X=-0.19 $Y=1.66 $X2=5.64 $Y2=1.585
cc_97 VPB N_A1_c_329_n 0.0490405f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.795
cc_98 VPB A1 0.00393152f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=2.46
cc_99 VPB N_A_31_94#_c_359_n 0.0453626f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=2.46
cc_100 VPB N_A_31_94#_c_361_n 0.0429428f $X=-0.19 $Y=1.66 $X2=3.015 $Y2=2.46
cc_101 VPB N_A_31_94#_c_369_n 0.0342569f $X=-0.19 $Y=1.66 $X2=1.655 $Y2=0.505
cc_102 VPB N_A_31_94#_c_370_n 0.0194882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_31_94#_c_371_n 0.00267616f $X=-0.19 $Y=1.66 $X2=3.105 $Y2=1.195
cc_104 VPB N_A_31_94#_c_372_n 0.0115102f $X=-0.19 $Y=1.66 $X2=5.61 $Y2=1.28
cc_105 VPB N_A_31_94#_c_373_n 0.00219628f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=1.195
cc_106 VPB N_A_31_94#_c_364_n 0.0100109f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.195
cc_107 VPB N_A_31_94#_c_365_n 0.00690382f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.385
cc_108 VPB N_A_31_94#_c_366_n 0.0130153f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.55
cc_109 VPB N_A0_c_482_n 0.0351947f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=2.46
cc_110 VPB A0 0.00181321f $X=-0.19 $Y=1.66 $X2=1.59 $Y2=0.74
cc_111 VPB N_A3_c_519_n 0.0422683f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.795
cc_112 VPB A3 0.0052366f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=2.46
cc_113 VPB N_A2_c_552_n 0.00730095f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.795
cc_114 VPB N_A2_c_557_n 0.0239954f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.885
cc_115 VPB A2 0.0041529f $X=-0.19 $Y=1.66 $X2=1.59 $Y2=1.26
cc_116 VPB N_A_1500_94#_c_601_n 0.0177252f $X=-0.19 $Y=1.66 $X2=1.59 $Y2=0.74
cc_117 VPB N_A_1500_94#_c_597_n 0.00852657f $X=-0.19 $Y=1.66 $X2=3.015 $Y2=2.46
cc_118 VPB N_A_1500_94#_c_603_n 0.00745992f $X=-0.19 $Y=1.66 $X2=1.57 $Y2=1.11
cc_119 VPB N_A_1500_94#_c_599_n 0.00134659f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=0.59
cc_120 VPB N_A_1500_94#_c_600_n 0.0278524f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=1.11
cc_121 VPB N_S1_c_651_n 0.0324895f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.795
cc_122 VPB N_S1_c_656_n 0.00664335f $X=-0.19 $Y=1.66 $X2=3.015 $Y2=2.46
cc_123 VPB N_S1_c_660_n 0.0267723f $X=-0.19 $Y=1.66 $X2=4.47 $Y2=1.22
cc_124 VPB S1 0.00543304f $X=-0.19 $Y=1.66 $X2=5.685 $Y2=2.46
cc_125 VPB N_A_1429_74#_c_736_n 0.0167473f $X=-0.19 $Y=1.66 $X2=1.59 $Y2=0.74
cc_126 VPB N_A_1429_74#_c_737_n 0.0176404f $X=-0.19 $Y=1.66 $X2=4.47 $Y2=1.22
cc_127 VPB N_A_1429_74#_c_730_n 0.0187083f $X=-0.19 $Y=1.66 $X2=5.685 $Y2=1.885
cc_128 VPB N_A_1429_74#_c_731_n 0.0167509f $X=-0.19 $Y=1.66 $X2=1.57 $Y2=0.59
cc_129 VPB N_A_1429_74#_c_740_n 0.0179765f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=0.59
cc_130 VPB N_A_1429_74#_c_741_n 0.00465423f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=1.615
cc_131 VPB N_A_1429_74#_c_742_n 0.00216079f $X=-0.19 $Y=1.66 $X2=5.61 $Y2=1.585
cc_132 VPB N_A_1429_74#_c_735_n 3.82886e-19 $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.425
cc_133 VPB N_VPWR_c_833_n 0.0154382f $X=-0.19 $Y=1.66 $X2=4.47 $Y2=0.74
cc_134 VPB N_VPWR_c_834_n 0.00990533f $X=-0.19 $Y=1.66 $X2=2.835 $Y2=0.505
cc_135 VPB N_VPWR_c_835_n 0.0113419f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=1.28
cc_136 VPB N_VPWR_c_836_n 0.0707244f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=1.615
cc_137 VPB N_VPWR_c_837_n 0.00808684f $X=-0.19 $Y=1.66 $X2=3.105 $Y2=1.195
cc_138 VPB N_VPWR_c_838_n 0.0104926f $X=-0.19 $Y=1.66 $X2=5.61 $Y2=1.585
cc_139 VPB N_VPWR_c_839_n 0.0595963f $X=-0.19 $Y=1.66 $X2=5.64 $Y2=1.585
cc_140 VPB N_VPWR_c_840_n 0.0236066f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.425
cc_141 VPB N_VPWR_c_841_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.425
cc_142 VPB N_VPWR_c_842_n 0.0730403f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.195
cc_143 VPB N_VPWR_c_843_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_844_n 0.0643736f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.425
cc_145 VPB N_VPWR_c_845_n 0.0204479f $X=-0.19 $Y=1.66 $X2=5.64 $Y2=1.585
cc_146 VPB N_VPWR_c_846_n 0.00614248f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.385
cc_147 VPB N_VPWR_c_847_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_832_n 0.168319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_333_74#_c_937_n 0.0067852f $X=-0.19 $Y=1.66 $X2=5.685 $Y2=1.885
cc_150 VPB N_A_333_74#_c_938_n 0.00452641f $X=-0.19 $Y=1.66 $X2=1.655 $Y2=0.505
cc_151 VPB N_A_333_74#_c_939_n 0.0020925f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=0.59
cc_152 VPB N_A_333_74#_c_933_n 0.00704428f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=1.28
cc_153 VPB N_A_333_74#_c_941_n 0.00382315f $X=-0.19 $Y=1.66 $X2=5.475 $Y2=1.195
cc_154 VPB N_A_333_74#_c_942_n 0.0164543f $X=-0.19 $Y=1.66 $X2=5.61 $Y2=1.28
cc_155 VPB N_A_333_74#_c_936_n 0.00506387f $X=-0.19 $Y=1.66 $X2=5.61 $Y2=1.585
cc_156 VPB N_A_333_74#_c_944_n 0.00326467f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.195
cc_157 VPB N_A_909_74#_c_1072_n 0.00843508f $X=-0.19 $Y=1.66 $X2=5.685 $Y2=1.885
cc_158 VPB N_A_909_74#_c_1073_n 0.0060908f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=1.615
cc_159 VPB N_A_909_74#_c_1074_n 0.0112726f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=1.615
cc_160 VPB N_A_909_74#_c_1068_n 0.00219993f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=1.195
cc_161 VPB N_A_909_74#_c_1076_n 0.00273342f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.195
cc_162 VPB X 5.28262e-19 $X=-0.19 $Y=1.66 $X2=0.645 $Y2=2.46
cc_163 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=1.195
cc_164 N_S0_M1010_g N_A1_M1013_g 0.0618951f $X=1.59 $Y=0.74 $X2=0 $Y2=0
cc_165 N_S0_c_173_n N_A1_M1013_g 0.0166126f $X=1.485 $Y=1.195 $X2=0 $Y2=0
cc_166 S0 N_A1_M1013_g 0.00165651f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_167 N_S0_c_179_n N_A1_M1013_g 0.00701358f $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_168 N_S0_c_180_n N_A1_M1013_g 0.00939458f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_169 N_S0_c_165_n N_A1_c_329_n 0.0155236f $X=0.645 $Y=1.795 $X2=0 $Y2=0
cc_170 N_S0_c_183_n N_A1_c_329_n 0.023133f $X=0.645 $Y=1.885 $X2=0 $Y2=0
cc_171 N_S0_c_173_n N_A1_c_329_n 0.0051813f $X=1.485 $Y=1.195 $X2=0 $Y2=0
cc_172 N_S0_c_174_n N_A1_c_329_n 0.0090888f $X=1.68 $Y=1.425 $X2=0 $Y2=0
cc_173 S0 N_A1_c_329_n 3.31425e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_174 N_S0_c_179_n N_A1_c_329_n 0.00649335f $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_175 N_S0_c_165_n A1 0.00150864f $X=0.645 $Y=1.795 $X2=0 $Y2=0
cc_176 N_S0_c_173_n A1 0.0368142f $X=1.485 $Y=1.195 $X2=0 $Y2=0
cc_177 N_S0_c_174_n A1 4.25896e-19 $X=1.68 $Y=1.425 $X2=0 $Y2=0
cc_178 S0 A1 0.00800143f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_179 N_S0_c_167_n N_A_31_94#_c_359_n 0.0318299f $X=3.015 $Y=1.885 $X2=0 $Y2=0
cc_180 N_S0_c_174_n N_A_31_94#_c_359_n 0.00910163f $X=1.68 $Y=1.425 $X2=0 $Y2=0
cc_181 N_S0_M1010_g N_A_31_94#_M1014_g 0.0153356f $X=1.59 $Y=0.74 $X2=0 $Y2=0
cc_182 N_S0_c_206_p N_A_31_94#_M1014_g 0.0137849f $X=2.835 $Y=0.505 $X2=0 $Y2=0
cc_183 N_S0_c_207_p N_A_31_94#_M1014_g 0.00721875f $X=2.97 $Y=1.11 $X2=0 $Y2=0
cc_184 N_S0_c_169_n N_A_31_94#_M1014_g 9.0572e-19 $X=2.94 $Y=1.615 $X2=0 $Y2=0
cc_185 N_S0_c_173_n N_A_31_94#_M1014_g 7.08885e-19 $X=1.485 $Y=1.195 $X2=0 $Y2=0
cc_186 N_S0_c_174_n N_A_31_94#_M1014_g 0.00322529f $X=1.68 $Y=1.425 $X2=0 $Y2=0
cc_187 N_S0_c_175_n N_A_31_94#_M1014_g 9.92616e-19 $X=2.97 $Y=1.195 $X2=0 $Y2=0
cc_188 N_S0_c_168_n N_A_31_94#_c_361_n 0.0440592f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_189 N_S0_c_171_n N_A_31_94#_c_361_n 0.00143877f $X=5.475 $Y=1.195 $X2=0 $Y2=0
cc_190 N_S0_c_172_n N_A_31_94#_c_361_n 0.00101098f $X=5.64 $Y=1.585 $X2=0 $Y2=0
cc_191 N_S0_c_177_n N_A_31_94#_c_361_n 0.00565283f $X=4.56 $Y=1.385 $X2=0 $Y2=0
cc_192 N_S0_c_168_n N_A_31_94#_M1005_g 0.00221213f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_193 N_S0_c_171_n N_A_31_94#_M1005_g 0.012897f $X=5.475 $Y=1.195 $X2=0 $Y2=0
cc_194 N_S0_c_172_n N_A_31_94#_M1005_g 0.00493866f $X=5.64 $Y=1.585 $X2=0 $Y2=0
cc_195 N_S0_c_176_n N_A_31_94#_M1005_g 0.00120505f $X=4.56 $Y=1.195 $X2=0 $Y2=0
cc_196 N_S0_c_177_n N_A_31_94#_M1005_g 0.00855265f $X=4.56 $Y=1.385 $X2=0 $Y2=0
cc_197 N_S0_c_181_n N_A_31_94#_M1005_g 0.0194574f $X=4.56 $Y=1.22 $X2=0 $Y2=0
cc_198 N_S0_c_183_n N_A_31_94#_c_369_n 0.00853629f $X=0.645 $Y=1.885 $X2=0 $Y2=0
cc_199 S0 N_A_31_94#_c_363_n 0.00211202f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_200 N_S0_c_180_n N_A_31_94#_c_363_n 0.0113051f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_201 N_S0_c_183_n N_A_31_94#_c_399_n 0.00892277f $X=0.645 $Y=1.885 $X2=0 $Y2=0
cc_202 N_S0_c_173_n N_A_31_94#_c_399_n 0.0136162f $X=1.485 $Y=1.195 $X2=0 $Y2=0
cc_203 S0 N_A_31_94#_c_399_n 0.00689942f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_204 N_S0_c_169_n N_A_31_94#_c_402_n 0.0021071f $X=2.94 $Y=1.615 $X2=0 $Y2=0
cc_205 N_S0_c_176_n N_A_31_94#_c_402_n 0.0117141f $X=4.56 $Y=1.195 $X2=0 $Y2=0
cc_206 N_S0_c_183_n N_A_31_94#_c_372_n 0.00381008f $X=0.645 $Y=1.885 $X2=0 $Y2=0
cc_207 S0 N_A_31_94#_c_372_n 0.00602207f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_208 N_S0_c_179_n N_A_31_94#_c_372_n 8.51315e-19 $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_209 N_S0_c_173_n N_A_31_94#_c_364_n 0.00978474f $X=1.485 $Y=1.195 $X2=0 $Y2=0
cc_210 N_S0_c_174_n N_A_31_94#_c_364_n 4.67042e-19 $X=1.68 $Y=1.425 $X2=0 $Y2=0
cc_211 N_S0_c_168_n N_A_31_94#_c_365_n 0.00482589f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_212 N_S0_c_171_n N_A_31_94#_c_365_n 0.0253679f $X=5.475 $Y=1.195 $X2=0 $Y2=0
cc_213 N_S0_c_172_n N_A_31_94#_c_365_n 0.0181422f $X=5.64 $Y=1.585 $X2=0 $Y2=0
cc_214 N_S0_c_176_n N_A_31_94#_c_365_n 0.00632157f $X=4.56 $Y=1.195 $X2=0 $Y2=0
cc_215 N_S0_c_177_n N_A_31_94#_c_365_n 5.14735e-19 $X=4.56 $Y=1.385 $X2=0 $Y2=0
cc_216 N_S0_c_165_n N_A_31_94#_c_366_n 0.00980729f $X=0.645 $Y=1.795 $X2=0 $Y2=0
cc_217 S0 N_A_31_94#_c_366_n 0.0321761f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_218 N_S0_c_179_n N_A_31_94#_c_366_n 0.00232633f $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_219 N_S0_c_180_n N_A_31_94#_c_366_n 0.00346005f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_220 N_S0_c_206_p N_A0_M1023_g 0.00365122f $X=2.835 $Y=0.505 $X2=0 $Y2=0
cc_221 N_S0_c_207_p N_A0_M1023_g 0.013009f $X=2.97 $Y=1.11 $X2=0 $Y2=0
cc_222 N_S0_c_170_n N_A0_M1023_g 0.0130662f $X=4.395 $Y=1.195 $X2=0 $Y2=0
cc_223 N_S0_c_169_n N_A0_c_480_n 0.00639658f $X=2.94 $Y=1.615 $X2=0 $Y2=0
cc_224 N_S0_c_170_n N_A0_c_480_n 0.0101907f $X=4.395 $Y=1.195 $X2=0 $Y2=0
cc_225 N_S0_c_167_n N_A0_c_481_n 0.0207461f $X=3.015 $Y=1.885 $X2=0 $Y2=0
cc_226 N_S0_c_169_n N_A0_c_481_n 4.14716e-19 $X=2.94 $Y=1.615 $X2=0 $Y2=0
cc_227 N_S0_c_167_n N_A0_c_482_n 0.063142f $X=3.015 $Y=1.885 $X2=0 $Y2=0
cc_228 N_S0_c_167_n A0 0.00114283f $X=3.015 $Y=1.885 $X2=0 $Y2=0
cc_229 N_S0_c_169_n A0 0.0207106f $X=2.94 $Y=1.615 $X2=0 $Y2=0
cc_230 N_S0_c_170_n A0 0.0267376f $X=4.395 $Y=1.195 $X2=0 $Y2=0
cc_231 N_S0_c_170_n N_A3_M1019_g 0.0156888f $X=4.395 $Y=1.195 $X2=0 $Y2=0
cc_232 N_S0_c_176_n N_A3_M1019_g 0.00121532f $X=4.56 $Y=1.195 $X2=0 $Y2=0
cc_233 N_S0_c_181_n N_A3_M1019_g 0.063939f $X=4.56 $Y=1.22 $X2=0 $Y2=0
cc_234 N_S0_c_170_n N_A3_c_519_n 0.00427011f $X=4.395 $Y=1.195 $X2=0 $Y2=0
cc_235 N_S0_c_177_n N_A3_c_519_n 0.0062914f $X=4.56 $Y=1.385 $X2=0 $Y2=0
cc_236 N_S0_c_170_n A3 0.0250329f $X=4.395 $Y=1.195 $X2=0 $Y2=0
cc_237 N_S0_c_176_n A3 0.00698305f $X=4.56 $Y=1.195 $X2=0 $Y2=0
cc_238 N_S0_c_177_n A3 5.6641e-19 $X=4.56 $Y=1.385 $X2=0 $Y2=0
cc_239 N_S0_c_168_n N_A2_c_552_n 0.00777699f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_240 N_S0_c_168_n N_A2_c_557_n 0.0539138f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_241 N_S0_c_168_n A2 0.0025277f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_242 N_S0_c_171_n A2 0.00901589f $X=5.475 $Y=1.195 $X2=0 $Y2=0
cc_243 N_S0_c_172_n A2 0.0379793f $X=5.64 $Y=1.585 $X2=0 $Y2=0
cc_244 N_S0_c_168_n N_A2_c_554_n 0.0203953f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_245 N_S0_c_172_n N_A2_c_554_n 0.00109924f $X=5.64 $Y=1.585 $X2=0 $Y2=0
cc_246 N_S0_c_171_n N_A2_c_555_n 0.00320079f $X=5.475 $Y=1.195 $X2=0 $Y2=0
cc_247 N_S0_c_183_n N_VPWR_c_833_n 0.0101886f $X=0.645 $Y=1.885 $X2=0 $Y2=0
cc_248 N_S0_c_173_n N_VPWR_c_833_n 0.00387653f $X=1.485 $Y=1.195 $X2=0 $Y2=0
cc_249 S0 N_VPWR_c_833_n 0.00199233f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_250 N_S0_c_168_n N_VPWR_c_835_n 8.81747e-19 $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_251 N_S0_c_183_n N_VPWR_c_840_n 0.00445602f $X=0.645 $Y=1.885 $X2=0 $Y2=0
cc_252 N_S0_c_167_n N_VPWR_c_842_n 0.00291513f $X=3.015 $Y=1.885 $X2=0 $Y2=0
cc_253 N_S0_c_168_n N_VPWR_c_844_n 0.00300876f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_254 N_S0_c_183_n N_VPWR_c_832_n 0.00862058f $X=0.645 $Y=1.885 $X2=0 $Y2=0
cc_255 N_S0_c_167_n N_VPWR_c_832_n 0.00361222f $X=3.015 $Y=1.885 $X2=0 $Y2=0
cc_256 N_S0_c_168_n N_VPWR_c_832_n 0.00370553f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_257 N_S0_c_206_p N_A_333_74#_M1010_d 0.0185809f $X=2.835 $Y=0.505 $X2=-0.19
+ $Y2=-0.245
cc_258 N_S0_M1010_g N_A_333_74#_c_946_n 0.00343798f $X=1.59 $Y=0.74 $X2=0 $Y2=0
cc_259 N_S0_c_283_p N_A_333_74#_c_946_n 0.0232888f $X=1.57 $Y=1.11 $X2=0 $Y2=0
cc_260 N_S0_c_206_p N_A_333_74#_c_946_n 0.0514462f $X=2.835 $Y=0.505 $X2=0 $Y2=0
cc_261 N_S0_c_207_p N_A_333_74#_c_946_n 0.0277115f $X=2.97 $Y=1.11 $X2=0 $Y2=0
cc_262 N_S0_c_170_n N_A_333_74#_c_937_n 0.00774188f $X=4.395 $Y=1.195 $X2=0
+ $Y2=0
cc_263 N_S0_c_168_n N_A_333_74#_c_938_n 0.0142816f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_264 N_S0_c_172_n N_A_333_74#_c_938_n 0.00895395f $X=5.64 $Y=1.585 $X2=0 $Y2=0
cc_265 N_S0_c_168_n N_A_333_74#_c_939_n 7.56472e-19 $X=5.685 $Y=1.885 $X2=0
+ $Y2=0
cc_266 N_S0_c_172_n N_A_333_74#_c_939_n 0.00738039f $X=5.64 $Y=1.585 $X2=0 $Y2=0
cc_267 N_S0_c_167_n N_A_333_74#_c_942_n 0.0519836f $X=3.015 $Y=1.885 $X2=0 $Y2=0
cc_268 N_S0_c_169_n N_A_333_74#_c_942_n 0.0211718f $X=2.94 $Y=1.615 $X2=0 $Y2=0
cc_269 N_S0_c_170_n N_A_333_74#_c_942_n 0.00676946f $X=4.395 $Y=1.195 $X2=0
+ $Y2=0
cc_270 N_S0_c_167_n N_A_333_74#_c_936_n 0.00599691f $X=3.015 $Y=1.885 $X2=0
+ $Y2=0
cc_271 N_S0_c_207_p N_A_333_74#_c_936_n 0.00142951f $X=2.97 $Y=1.11 $X2=0 $Y2=0
cc_272 N_S0_c_169_n N_A_333_74#_c_936_n 0.0376502f $X=2.94 $Y=1.615 $X2=0 $Y2=0
cc_273 N_S0_c_173_n N_A_333_74#_c_936_n 0.00449018f $X=1.485 $Y=1.195 $X2=0
+ $Y2=0
cc_274 N_S0_c_174_n N_A_333_74#_c_936_n 2.08099e-19 $X=1.68 $Y=1.425 $X2=0 $Y2=0
cc_275 N_S0_c_175_n N_A_333_74#_c_936_n 0.0143571f $X=2.97 $Y=1.195 $X2=0 $Y2=0
cc_276 N_S0_c_176_n N_A_909_74#_M1016_d 0.00195473f $X=4.56 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_277 N_S0_c_168_n N_A_909_74#_c_1078_n 0.0144091f $X=5.685 $Y=1.885 $X2=0
+ $Y2=0
cc_278 N_S0_c_168_n N_A_909_74#_c_1065_n 0.00266197f $X=5.685 $Y=1.885 $X2=0
+ $Y2=0
cc_279 N_S0_c_171_n N_A_909_74#_c_1065_n 0.046315f $X=5.475 $Y=1.195 $X2=0 $Y2=0
cc_280 N_S0_c_171_n N_A_909_74#_c_1069_n 0.0283569f $X=5.475 $Y=1.195 $X2=0
+ $Y2=0
cc_281 N_S0_c_176_n N_A_909_74#_c_1069_n 0.0140846f $X=4.56 $Y=1.195 $X2=0 $Y2=0
cc_282 N_S0_c_177_n N_A_909_74#_c_1069_n 9.23826e-19 $X=4.56 $Y=1.385 $X2=0
+ $Y2=0
cc_283 N_S0_c_181_n N_A_909_74#_c_1069_n 0.0216345f $X=4.56 $Y=1.22 $X2=0 $Y2=0
cc_284 S0 N_VGND_M1001_d 0.00727922f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_285 N_S0_M1010_g N_VGND_c_1222_n 0.00144364f $X=1.59 $Y=0.74 $X2=0 $Y2=0
cc_286 N_S0_c_173_n N_VGND_c_1222_n 0.0246662f $X=1.485 $Y=1.195 $X2=0 $Y2=0
cc_287 N_S0_c_180_n N_VGND_c_1222_n 0.00808843f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_288 N_S0_c_206_p N_VGND_c_1223_n 0.00845662f $X=2.835 $Y=0.505 $X2=0 $Y2=0
cc_289 N_S0_c_207_p N_VGND_c_1223_n 0.0161363f $X=2.97 $Y=1.11 $X2=0 $Y2=0
cc_290 N_S0_c_170_n N_VGND_c_1223_n 0.0368014f $X=4.395 $Y=1.195 $X2=0 $Y2=0
cc_291 N_S0_c_180_n N_VGND_c_1228_n 0.00486269f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_292 N_S0_c_181_n N_VGND_c_1230_n 0.00445602f $X=4.56 $Y=1.22 $X2=0 $Y2=0
cc_293 N_S0_M1010_g N_VGND_c_1232_n 0.00300757f $X=1.59 $Y=0.74 $X2=0 $Y2=0
cc_294 N_S0_c_206_p N_VGND_c_1232_n 0.0428549f $X=2.835 $Y=0.505 $X2=0 $Y2=0
cc_295 N_S0_c_319_p N_VGND_c_1232_n 0.00503142f $X=1.655 $Y=0.505 $X2=0 $Y2=0
cc_296 N_S0_M1010_g N_VGND_c_1237_n 0.00371003f $X=1.59 $Y=0.74 $X2=0 $Y2=0
cc_297 N_S0_c_206_p N_VGND_c_1237_n 0.0484519f $X=2.835 $Y=0.505 $X2=0 $Y2=0
cc_298 N_S0_c_319_p N_VGND_c_1237_n 0.00531343f $X=1.655 $Y=0.505 $X2=0 $Y2=0
cc_299 N_S0_c_180_n N_VGND_c_1237_n 0.00514438f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_300 N_S0_c_181_n N_VGND_c_1237_n 0.008597f $X=4.56 $Y=1.22 $X2=0 $Y2=0
cc_301 N_S0_c_206_p A_507_74# 0.0196082f $X=2.835 $Y=0.505 $X2=-0.19 $Y2=-0.245
cc_302 N_S0_c_207_p A_507_74# 0.0192269f $X=2.97 $Y=1.11 $X2=-0.19 $Y2=-0.245
cc_303 N_S0_c_171_n A_1047_74# 0.00296756f $X=5.475 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_304 N_A1_c_329_n N_A_31_94#_c_359_n 8.28942e-19 $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_305 N_A1_c_329_n N_A_31_94#_c_399_n 0.0145894f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_306 A1 N_A_31_94#_c_399_n 0.010433f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_307 N_A1_c_329_n N_A_31_94#_c_372_n 3.53657e-19 $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_308 N_A1_c_329_n N_VPWR_c_833_n 0.0337103f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_309 A1 N_VPWR_c_833_n 0.00844532f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_310 N_A1_c_329_n N_VPWR_c_842_n 0.00461464f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_311 N_A1_c_329_n N_VPWR_c_832_n 0.00915467f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_312 N_A1_M1013_g N_VGND_c_1222_n 0.0135991f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A1_M1013_g N_VGND_c_1232_n 0.00383152f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A1_M1013_g N_VGND_c_1237_n 0.0075725f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A_31_94#_c_402_n A0 0.00274892f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_316 N_A_31_94#_c_361_n N_A3_c_519_n 0.0215292f $X=4.995 $Y=1.885 $X2=0 $Y2=0
cc_317 N_A_31_94#_c_402_n A3 0.00251567f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_318 N_A_31_94#_M1005_g A2 4.44262e-19 $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A_31_94#_c_365_n A2 8.70553e-19 $X=5.1 $Y=1.625 $X2=0 $Y2=0
cc_320 N_A_31_94#_c_399_n N_VPWR_M1007_d 0.00561589f $X=2.015 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_321 N_A_31_94#_c_399_n N_VPWR_c_833_n 0.0375103f $X=2.015 $Y=2.035 $X2=0
+ $Y2=0
cc_322 N_A_31_94#_c_370_n N_VPWR_c_833_n 3.02414e-19 $X=0.385 $Y=2.035 $X2=0
+ $Y2=0
cc_323 N_A_31_94#_c_372_n N_VPWR_c_833_n 0.0417249f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_324 N_A_31_94#_c_402_n N_VPWR_c_834_n 0.0027508f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_325 N_A_31_94#_c_369_n N_VPWR_c_840_n 0.0145938f $X=0.42 $Y=2.815 $X2=0 $Y2=0
cc_326 N_A_31_94#_c_359_n N_VPWR_c_842_n 0.00461464f $X=2.295 $Y=1.885 $X2=0
+ $Y2=0
cc_327 N_A_31_94#_c_361_n N_VPWR_c_844_n 0.00445405f $X=4.995 $Y=1.885 $X2=0
+ $Y2=0
cc_328 N_A_31_94#_c_359_n N_VPWR_c_832_n 0.0091652f $X=2.295 $Y=1.885 $X2=0
+ $Y2=0
cc_329 N_A_31_94#_c_361_n N_VPWR_c_832_n 0.0045994f $X=4.995 $Y=1.885 $X2=0
+ $Y2=0
cc_330 N_A_31_94#_c_369_n N_VPWR_c_832_n 0.0120466f $X=0.42 $Y=2.815 $X2=0 $Y2=0
cc_331 N_A_31_94#_c_399_n A_264_392# 0.0445093f $X=2.015 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_332 N_A_31_94#_c_371_n A_264_392# 0.00793794f $X=2.305 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_333 N_A_31_94#_c_364_n A_264_392# 0.00524585f $X=2.22 $Y=1.615 $X2=-0.19
+ $Y2=-0.245
cc_334 N_A_31_94#_c_402_n N_A_333_74#_M1000_d 0.00687888f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_335 N_A_31_94#_c_359_n N_A_333_74#_c_946_n 0.00297754f $X=2.295 $Y=1.885
+ $X2=0 $Y2=0
cc_336 N_A_31_94#_M1014_g N_A_333_74#_c_946_n 0.023686f $X=2.46 $Y=0.74 $X2=0
+ $Y2=0
cc_337 N_A_31_94#_c_364_n N_A_333_74#_c_946_n 0.0129016f $X=2.22 $Y=1.615 $X2=0
+ $Y2=0
cc_338 N_A_31_94#_c_361_n N_A_333_74#_c_937_n 7.52993e-19 $X=4.995 $Y=1.885
+ $X2=0 $Y2=0
cc_339 N_A_31_94#_c_402_n N_A_333_74#_c_937_n 0.0598959f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_340 N_A_31_94#_c_373_n N_A_333_74#_c_937_n 6.89416e-19 $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_341 N_A_31_94#_c_365_n N_A_333_74#_c_937_n 0.00200875f $X=5.1 $Y=1.625 $X2=0
+ $Y2=0
cc_342 N_A_31_94#_c_361_n N_A_333_74#_c_972_n 0.00253283f $X=4.995 $Y=1.885
+ $X2=0 $Y2=0
cc_343 N_A_31_94#_c_373_n N_A_333_74#_c_972_n 6.41773e-19 $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_344 N_A_31_94#_c_365_n N_A_333_74#_c_972_n 3.57346e-19 $X=5.1 $Y=1.625 $X2=0
+ $Y2=0
cc_345 N_A_31_94#_c_361_n N_A_333_74#_c_975_n 0.0144128f $X=4.995 $Y=1.885 $X2=0
+ $Y2=0
cc_346 N_A_31_94#_c_402_n N_A_333_74#_c_975_n 0.0264387f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_347 N_A_31_94#_c_373_n N_A_333_74#_c_975_n 0.00334834f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_348 N_A_31_94#_c_365_n N_A_333_74#_c_975_n 0.0200153f $X=5.1 $Y=1.625 $X2=0
+ $Y2=0
cc_349 N_A_31_94#_c_361_n N_A_333_74#_c_939_n 0.0037267f $X=4.995 $Y=1.885 $X2=0
+ $Y2=0
cc_350 N_A_31_94#_c_373_n N_A_333_74#_c_939_n 0.00113398f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_351 N_A_31_94#_c_365_n N_A_333_74#_c_939_n 0.0134674f $X=5.1 $Y=1.625 $X2=0
+ $Y2=0
cc_352 N_A_31_94#_c_402_n N_A_333_74#_c_942_n 0.0940841f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_353 N_A_31_94#_c_371_n N_A_333_74#_c_942_n 3.61668e-19 $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_354 N_A_31_94#_c_359_n N_A_333_74#_c_936_n 0.0357651f $X=2.295 $Y=1.885 $X2=0
+ $Y2=0
cc_355 N_A_31_94#_M1014_g N_A_333_74#_c_936_n 0.0171633f $X=2.46 $Y=0.74 $X2=0
+ $Y2=0
cc_356 N_A_31_94#_c_371_n N_A_333_74#_c_936_n 3.32471e-19 $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_357 N_A_31_94#_c_364_n N_A_333_74#_c_936_n 0.0501859f $X=2.22 $Y=1.615 $X2=0
+ $Y2=0
cc_358 N_A_31_94#_c_402_n A_840_392# 0.0212324f $X=4.895 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_359 N_A_31_94#_c_373_n A_840_392# 9.15431e-19 $X=5.04 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_360 N_A_31_94#_c_373_n N_A_909_74#_M1015_d 4.80017e-19 $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_361 N_A_31_94#_c_365_n N_A_909_74#_M1015_d 0.00294616f $X=5.1 $Y=1.625 $X2=0
+ $Y2=0
cc_362 N_A_31_94#_c_361_n N_A_909_74#_c_1078_n 0.0165226f $X=4.995 $Y=1.885
+ $X2=0 $Y2=0
cc_363 N_A_31_94#_M1005_g N_A_909_74#_c_1065_n 0.0111936f $X=5.16 $Y=0.74 $X2=0
+ $Y2=0
cc_364 N_A_31_94#_M1005_g N_A_909_74#_c_1069_n 0.0313844f $X=5.16 $Y=0.74 $X2=0
+ $Y2=0
cc_365 N_A_31_94#_c_363_n N_VGND_c_1222_n 0.0195703f $X=0.3 $Y=0.75 $X2=0 $Y2=0
cc_366 N_A_31_94#_c_363_n N_VGND_c_1228_n 0.00904149f $X=0.3 $Y=0.75 $X2=0 $Y2=0
cc_367 N_A_31_94#_M1005_g N_VGND_c_1230_n 0.00439937f $X=5.16 $Y=0.74 $X2=0
+ $Y2=0
cc_368 N_A_31_94#_M1014_g N_VGND_c_1232_n 0.00300876f $X=2.46 $Y=0.74 $X2=0
+ $Y2=0
cc_369 N_A_31_94#_M1014_g N_VGND_c_1237_n 0.00376442f $X=2.46 $Y=0.74 $X2=0
+ $Y2=0
cc_370 N_A_31_94#_M1005_g N_VGND_c_1237_n 0.00441434f $X=5.16 $Y=0.74 $X2=0
+ $Y2=0
cc_371 N_A_31_94#_c_363_n N_VGND_c_1237_n 0.0122078f $X=0.3 $Y=0.75 $X2=0 $Y2=0
cc_372 N_A0_M1023_g N_A3_M1019_g 0.010938f $X=3.39 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A0_c_480_n N_A3_M1019_g 0.00857915f $X=3.48 $Y=1.405 $X2=0 $Y2=0
cc_374 N_A0_c_481_n N_A3_c_519_n 0.0213989f $X=3.48 $Y=1.615 $X2=0 $Y2=0
cc_375 N_A0_c_482_n N_A3_c_519_n 0.0211556f $X=3.435 $Y=1.885 $X2=0 $Y2=0
cc_376 A0 N_A3_c_519_n 0.00109805f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_377 N_A0_c_481_n A3 3.7716e-19 $X=3.48 $Y=1.615 $X2=0 $Y2=0
cc_378 A0 A3 0.0265098f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_379 N_A0_c_482_n N_VPWR_c_834_n 0.0096544f $X=3.435 $Y=1.885 $X2=0 $Y2=0
cc_380 N_A0_c_482_n N_VPWR_c_842_n 0.00366292f $X=3.435 $Y=1.885 $X2=0 $Y2=0
cc_381 N_A0_c_482_n N_VPWR_c_832_n 0.00603185f $X=3.435 $Y=1.885 $X2=0 $Y2=0
cc_382 N_A0_c_482_n N_A_333_74#_c_937_n 0.0113712f $X=3.435 $Y=1.885 $X2=0 $Y2=0
cc_383 A0 N_A_333_74#_c_937_n 0.0162757f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_384 N_A0_c_482_n N_A_333_74#_c_972_n 5.78365e-19 $X=3.435 $Y=1.885 $X2=0
+ $Y2=0
cc_385 N_A0_c_482_n N_A_333_74#_c_942_n 0.0306844f $X=3.435 $Y=1.885 $X2=0 $Y2=0
cc_386 A0 N_A_333_74#_c_942_n 0.00961603f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_387 N_A0_M1023_g N_A_333_74#_c_936_n 4.86218e-19 $X=3.39 $Y=0.74 $X2=0 $Y2=0
cc_388 N_A0_M1023_g N_VGND_c_1223_n 0.0184517f $X=3.39 $Y=0.74 $X2=0 $Y2=0
cc_389 N_A0_c_480_n N_VGND_c_1223_n 8.94887e-19 $X=3.48 $Y=1.405 $X2=0 $Y2=0
cc_390 N_A0_M1023_g N_VGND_c_1232_n 0.00398535f $X=3.39 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A0_M1023_g N_VGND_c_1237_n 0.00792533f $X=3.39 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A3_c_519_n N_VPWR_c_834_n 0.0188446f $X=4.125 $Y=1.885 $X2=0 $Y2=0
cc_393 N_A3_c_519_n N_VPWR_c_844_n 0.00461464f $X=4.125 $Y=1.885 $X2=0 $Y2=0
cc_394 N_A3_c_519_n N_VPWR_c_832_n 0.00662122f $X=4.125 $Y=1.885 $X2=0 $Y2=0
cc_395 N_A3_c_519_n N_A_333_74#_c_937_n 0.0170944f $X=4.125 $Y=1.885 $X2=0 $Y2=0
cc_396 A3 N_A_333_74#_c_937_n 0.0232272f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_397 N_A3_c_519_n N_A_333_74#_c_972_n 0.00712777f $X=4.125 $Y=1.885 $X2=0
+ $Y2=0
cc_398 N_A3_c_519_n N_A_333_74#_c_997_n 0.00825839f $X=4.125 $Y=1.885 $X2=0
+ $Y2=0
cc_399 N_A3_c_519_n N_A_333_74#_c_942_n 7.7688e-19 $X=4.125 $Y=1.885 $X2=0 $Y2=0
cc_400 N_A3_M1019_g N_A_909_74#_c_1069_n 0.0017175f $X=4.08 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A3_M1019_g N_VGND_c_1223_n 0.0133278f $X=4.08 $Y=0.74 $X2=0 $Y2=0
cc_402 N_A3_M1019_g N_VGND_c_1230_n 0.00461464f $X=4.08 $Y=0.74 $X2=0 $Y2=0
cc_403 N_A3_M1019_g N_VGND_c_1237_n 0.00910635f $X=4.08 $Y=0.74 $X2=0 $Y2=0
cc_404 A2 N_S1_M1009_g 2.08945e-19 $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_405 N_A2_c_554_n N_S1_M1009_g 0.00250766f $X=6.18 $Y=1.385 $X2=0 $Y2=0
cc_406 N_A2_c_552_n N_S1_c_651_n 0.00219236f $X=6.105 $Y=1.795 $X2=0 $Y2=0
cc_407 N_A2_c_554_n N_S1_c_651_n 0.00153857f $X=6.18 $Y=1.385 $X2=0 $Y2=0
cc_408 N_A2_c_557_n N_VPWR_c_835_n 0.00835652f $X=6.105 $Y=1.885 $X2=0 $Y2=0
cc_409 N_A2_c_557_n N_VPWR_c_844_n 0.00413917f $X=6.105 $Y=1.885 $X2=0 $Y2=0
cc_410 N_A2_c_557_n N_VPWR_c_832_n 0.00402987f $X=6.105 $Y=1.885 $X2=0 $Y2=0
cc_411 N_A2_c_557_n N_A_333_74#_c_938_n 0.0160115f $X=6.105 $Y=1.885 $X2=0 $Y2=0
cc_412 A2 N_A_333_74#_c_938_n 0.0291858f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_413 N_A2_c_554_n N_A_333_74#_c_938_n 5.70384e-19 $X=6.18 $Y=1.385 $X2=0 $Y2=0
cc_414 N_A2_c_552_n N_A_333_74#_c_933_n 0.00365697f $X=6.105 $Y=1.795 $X2=0
+ $Y2=0
cc_415 N_A2_c_557_n N_A_333_74#_c_933_n 0.00175363f $X=6.105 $Y=1.885 $X2=0
+ $Y2=0
cc_416 A2 N_A_333_74#_c_933_n 0.0331323f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_417 N_A2_c_554_n N_A_333_74#_c_933_n 0.00259704f $X=6.18 $Y=1.385 $X2=0 $Y2=0
cc_418 A2 N_A_333_74#_c_934_n 0.00737832f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_419 N_A2_c_554_n N_A_333_74#_c_934_n 6.56322e-19 $X=6.18 $Y=1.385 $X2=0 $Y2=0
cc_420 N_A2_c_555_n N_A_333_74#_c_934_n 0.00247686f $X=6.18 $Y=1.22 $X2=0 $Y2=0
cc_421 N_A2_c_557_n N_A_333_74#_c_944_n 3.16517e-19 $X=6.105 $Y=1.885 $X2=0
+ $Y2=0
cc_422 A2 N_A_909_74#_c_1065_n 0.0231978f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_423 N_A2_c_554_n N_A_909_74#_c_1065_n 9.30761e-19 $X=6.18 $Y=1.385 $X2=0
+ $Y2=0
cc_424 N_A2_c_555_n N_A_909_74#_c_1065_n 0.0159612f $X=6.18 $Y=1.22 $X2=0 $Y2=0
cc_425 N_A2_c_557_n N_A_909_74#_c_1072_n 0.0125557f $X=6.105 $Y=1.885 $X2=0
+ $Y2=0
cc_426 N_A2_c_555_n N_A_909_74#_c_1066_n 0.0033505f $X=6.18 $Y=1.22 $X2=0 $Y2=0
cc_427 N_A2_c_557_n N_A_909_74#_c_1096_n 0.00558689f $X=6.105 $Y=1.885 $X2=0
+ $Y2=0
cc_428 N_A2_c_555_n N_VGND_c_1224_n 0.0189351f $X=6.18 $Y=1.22 $X2=0 $Y2=0
cc_429 N_A2_c_555_n N_VGND_c_1230_n 0.00383152f $X=6.18 $Y=1.22 $X2=0 $Y2=0
cc_430 N_A2_c_555_n N_VGND_c_1237_n 0.00374269f $X=6.18 $Y=1.22 $X2=0 $Y2=0
cc_431 N_A_1500_94#_c_596_n N_S1_M1009_g 0.0306434f $X=7.575 $Y=1.45 $X2=0 $Y2=0
cc_432 N_A_1500_94#_c_601_n N_S1_c_651_n 0.0352125f $X=7.59 $Y=1.885 $X2=0 $Y2=0
cc_433 N_A_1500_94#_c_597_n N_S1_c_651_n 0.0214393f $X=7.59 $Y=1.667 $X2=0 $Y2=0
cc_434 N_A_1500_94#_c_596_n N_S1_c_652_n 0.00976538f $X=7.575 $Y=1.45 $X2=0
+ $Y2=0
cc_435 N_A_1500_94#_c_598_n N_S1_M1008_g 0.00363246f $X=8.355 $Y=1.1 $X2=0 $Y2=0
cc_436 N_A_1500_94#_c_599_n N_S1_c_656_n 0.00123967f $X=8.23 $Y=1.615 $X2=0
+ $Y2=0
cc_437 N_A_1500_94#_c_600_n N_S1_c_656_n 0.0181406f $X=8.23 $Y=1.615 $X2=0 $Y2=0
cc_438 N_A_1500_94#_c_603_n N_S1_c_660_n 0.00417647f $X=8.365 $Y=2.155 $X2=0
+ $Y2=0
cc_439 N_A_1500_94#_c_597_n S1 0.0123956f $X=7.59 $Y=1.667 $X2=0 $Y2=0
cc_440 N_A_1500_94#_c_599_n S1 0.0276866f $X=8.23 $Y=1.615 $X2=0 $Y2=0
cc_441 N_A_1500_94#_c_596_n N_A_1429_74#_c_732_n 0.00150915f $X=7.575 $Y=1.45
+ $X2=0 $Y2=0
cc_442 N_A_1500_94#_M1018_s N_A_1429_74#_c_740_n 0.00438252f $X=8.225 $Y=1.94
+ $X2=0 $Y2=0
cc_443 N_A_1500_94#_c_601_n N_A_1429_74#_c_740_n 0.0101611f $X=7.59 $Y=1.885
+ $X2=0 $Y2=0
cc_444 N_A_1500_94#_c_596_n N_A_1429_74#_c_734_n 0.00359126f $X=7.575 $Y=1.45
+ $X2=0 $Y2=0
cc_445 N_A_1500_94#_c_601_n N_A_1429_74#_c_742_n 0.0100005f $X=7.59 $Y=1.885
+ $X2=0 $Y2=0
cc_446 N_A_1500_94#_c_601_n N_VPWR_c_836_n 0.00279479f $X=7.59 $Y=1.885 $X2=0
+ $Y2=0
cc_447 N_A_1500_94#_c_601_n N_VPWR_c_832_n 0.00357798f $X=7.59 $Y=1.885 $X2=0
+ $Y2=0
cc_448 N_A_1500_94#_c_596_n N_A_333_74#_c_935_n 0.0116708f $X=7.575 $Y=1.45
+ $X2=0 $Y2=0
cc_449 N_A_1500_94#_c_597_n N_A_333_74#_c_935_n 0.00686032f $X=7.59 $Y=1.667
+ $X2=0 $Y2=0
cc_450 N_A_1500_94#_c_598_n N_A_333_74#_c_935_n 0.0118332f $X=8.355 $Y=1.1 $X2=0
+ $Y2=0
cc_451 N_A_1500_94#_c_599_n N_A_333_74#_c_935_n 0.017009f $X=8.23 $Y=1.615 $X2=0
+ $Y2=0
cc_452 N_A_1500_94#_c_601_n N_A_333_74#_c_941_n 7.29978e-19 $X=7.59 $Y=1.885
+ $X2=0 $Y2=0
cc_453 N_A_1500_94#_c_601_n N_A_909_74#_c_1072_n 0.0120726f $X=7.59 $Y=1.885
+ $X2=0 $Y2=0
cc_454 N_A_1500_94#_c_596_n N_A_909_74#_c_1098_n 0.0121614f $X=7.575 $Y=1.45
+ $X2=0 $Y2=0
cc_455 N_A_1500_94#_c_601_n N_A_909_74#_c_1073_n 0.00791727f $X=7.59 $Y=1.885
+ $X2=0 $Y2=0
cc_456 N_A_1500_94#_c_597_n N_A_909_74#_c_1073_n 5.35718e-19 $X=7.59 $Y=1.667
+ $X2=0 $Y2=0
cc_457 N_A_1500_94#_c_603_n N_A_909_74#_c_1073_n 0.0285654f $X=8.365 $Y=2.155
+ $X2=0 $Y2=0
cc_458 N_A_1500_94#_c_599_n N_A_909_74#_c_1073_n 0.0213369f $X=8.23 $Y=1.615
+ $X2=0 $Y2=0
cc_459 N_A_1500_94#_c_600_n N_A_909_74#_c_1073_n 0.00722344f $X=8.23 $Y=1.615
+ $X2=0 $Y2=0
cc_460 N_A_1500_94#_M1018_s N_A_909_74#_c_1074_n 0.0138915f $X=8.225 $Y=1.94
+ $X2=0 $Y2=0
cc_461 N_A_1500_94#_c_603_n N_A_909_74#_c_1074_n 0.0202514f $X=8.365 $Y=2.155
+ $X2=0 $Y2=0
cc_462 N_A_1500_94#_M1008_s N_A_909_74#_c_1067_n 0.00964868f $X=8.205 $Y=0.6
+ $X2=0 $Y2=0
cc_463 N_A_1500_94#_c_598_n N_A_909_74#_c_1067_n 0.0214562f $X=8.355 $Y=1.1
+ $X2=0 $Y2=0
cc_464 N_A_1500_94#_c_600_n N_A_909_74#_c_1067_n 0.00429515f $X=8.23 $Y=1.615
+ $X2=0 $Y2=0
cc_465 N_A_1500_94#_c_598_n N_A_909_74#_c_1068_n 0.0281134f $X=8.355 $Y=1.1
+ $X2=0 $Y2=0
cc_466 N_A_1500_94#_c_603_n N_A_909_74#_c_1068_n 0.0298376f $X=8.365 $Y=2.155
+ $X2=0 $Y2=0
cc_467 N_A_1500_94#_c_599_n N_A_909_74#_c_1068_n 0.0278624f $X=8.23 $Y=1.615
+ $X2=0 $Y2=0
cc_468 N_A_1500_94#_c_600_n N_A_909_74#_c_1068_n 8.64189e-19 $X=8.23 $Y=1.615
+ $X2=0 $Y2=0
cc_469 N_A_1500_94#_c_601_n N_A_909_74#_c_1076_n 0.006161f $X=7.59 $Y=1.885
+ $X2=0 $Y2=0
cc_470 N_A_1500_94#_c_603_n N_A_909_74#_c_1076_n 0.00180878f $X=8.365 $Y=2.155
+ $X2=0 $Y2=0
cc_471 N_A_1500_94#_c_596_n N_A_909_74#_c_1071_n 0.00657413f $X=7.575 $Y=1.45
+ $X2=0 $Y2=0
cc_472 N_A_1500_94#_c_598_n N_A_909_74#_c_1071_n 3.89627e-19 $X=8.355 $Y=1.1
+ $X2=0 $Y2=0
cc_473 N_A_1500_94#_c_599_n N_A_909_74#_c_1071_n 0.00206203f $X=8.23 $Y=1.615
+ $X2=0 $Y2=0
cc_474 N_A_1500_94#_c_600_n N_A_909_74#_c_1071_n 0.0012069f $X=8.23 $Y=1.615
+ $X2=0 $Y2=0
cc_475 N_S1_c_655_n N_A_1429_74#_c_728_n 3.14814e-19 $X=8.725 $Y=1.405 $X2=0
+ $Y2=0
cc_476 N_S1_c_656_n N_A_1429_74#_c_736_n 7.65119e-19 $X=8.725 $Y=1.775 $X2=0
+ $Y2=0
cc_477 N_S1_c_655_n N_A_1429_74#_c_730_n 0.016675f $X=8.725 $Y=1.405 $X2=0 $Y2=0
cc_478 N_S1_c_656_n N_A_1429_74#_c_731_n 7.96211e-19 $X=8.725 $Y=1.775 $X2=0
+ $Y2=0
cc_479 N_S1_M1009_g N_A_1429_74#_c_732_n 3.76109e-19 $X=7.07 $Y=0.74 $X2=0 $Y2=0
cc_480 N_S1_c_652_n N_A_1429_74#_c_732_n 0.0293885f $X=8.635 $Y=0.185 $X2=0
+ $Y2=0
cc_481 N_S1_M1008_g N_A_1429_74#_c_732_n 0.0116641f $X=8.71 $Y=0.92 $X2=0 $Y2=0
cc_482 N_S1_c_660_n N_A_1429_74#_c_740_n 0.0140549f $X=8.725 $Y=1.865 $X2=0
+ $Y2=0
cc_483 N_S1_M1008_g N_A_1429_74#_c_733_n 0.010855f $X=8.71 $Y=0.92 $X2=0 $Y2=0
cc_484 N_S1_c_655_n N_A_1429_74#_c_733_n 3.56796e-19 $X=8.725 $Y=1.405 $X2=0
+ $Y2=0
cc_485 N_S1_c_656_n N_A_1429_74#_c_741_n 0.00188264f $X=8.725 $Y=1.775 $X2=0
+ $Y2=0
cc_486 N_S1_c_660_n N_A_1429_74#_c_741_n 0.0226543f $X=8.725 $Y=1.865 $X2=0
+ $Y2=0
cc_487 N_S1_M1009_g N_A_1429_74#_c_734_n 0.00719636f $X=7.07 $Y=0.74 $X2=0 $Y2=0
cc_488 N_S1_c_652_n N_A_1429_74#_c_734_n 0.00713661f $X=8.635 $Y=0.185 $X2=0
+ $Y2=0
cc_489 N_S1_c_653_n N_A_1429_74#_c_734_n 3.0179e-19 $X=7.145 $Y=0.185 $X2=0
+ $Y2=0
cc_490 N_S1_c_651_n N_A_1429_74#_c_742_n 0.017182f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_491 N_S1_c_655_n N_A_1429_74#_c_735_n 0.00197496f $X=8.725 $Y=1.405 $X2=0
+ $Y2=0
cc_492 N_S1_c_651_n N_VPWR_c_835_n 0.0092421f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_493 N_S1_c_651_n N_VPWR_c_836_n 0.00444353f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_494 N_S1_c_660_n N_VPWR_c_836_n 9.59479e-19 $X=8.725 $Y=1.865 $X2=0 $Y2=0
cc_495 N_S1_c_660_n N_VPWR_c_837_n 0.00182938f $X=8.725 $Y=1.865 $X2=0 $Y2=0
cc_496 N_S1_c_651_n N_VPWR_c_832_n 0.00448168f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_497 N_S1_M1009_g N_A_333_74#_c_933_n 0.00361032f $X=7.07 $Y=0.74 $X2=0 $Y2=0
cc_498 N_S1_c_651_n N_A_333_74#_c_933_n 0.00632618f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_499 S1 N_A_333_74#_c_933_n 0.0261339f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_500 N_S1_M1009_g N_A_333_74#_c_935_n 0.0122997f $X=7.07 $Y=0.74 $X2=0 $Y2=0
cc_501 N_S1_c_651_n N_A_333_74#_c_935_n 0.00433123f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_502 S1 N_A_333_74#_c_935_n 0.0471713f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_503 N_S1_c_651_n N_A_333_74#_c_941_n 0.00900412f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_504 S1 N_A_333_74#_c_941_n 0.0138774f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_505 N_S1_c_651_n N_A_909_74#_c_1072_n 0.0155288f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_506 S1 N_A_909_74#_c_1072_n 0.0122779f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_507 N_S1_M1009_g N_A_909_74#_c_1066_n 4.43891e-19 $X=7.07 $Y=0.74 $X2=0 $Y2=0
cc_508 N_S1_M1009_g N_A_909_74#_c_1098_n 0.00982569f $X=7.07 $Y=0.74 $X2=0 $Y2=0
cc_509 N_S1_c_652_n N_A_909_74#_c_1098_n 0.00159044f $X=8.635 $Y=0.185 $X2=0
+ $Y2=0
cc_510 N_S1_c_651_n N_A_909_74#_c_1073_n 0.0015462f $X=7.14 $Y=1.885 $X2=0 $Y2=0
cc_511 N_S1_c_660_n N_A_909_74#_c_1074_n 0.00917871f $X=8.725 $Y=1.865 $X2=0
+ $Y2=0
cc_512 N_S1_c_652_n N_A_909_74#_c_1067_n 0.00254292f $X=8.635 $Y=0.185 $X2=0
+ $Y2=0
cc_513 N_S1_M1008_g N_A_909_74#_c_1067_n 0.0107019f $X=8.71 $Y=0.92 $X2=0 $Y2=0
cc_514 N_S1_M1008_g N_A_909_74#_c_1068_n 0.023043f $X=8.71 $Y=0.92 $X2=0 $Y2=0
cc_515 N_S1_c_655_n N_A_909_74#_c_1068_n 0.00304199f $X=8.725 $Y=1.405 $X2=0
+ $Y2=0
cc_516 N_S1_c_656_n N_A_909_74#_c_1068_n 0.00862276f $X=8.725 $Y=1.775 $X2=0
+ $Y2=0
cc_517 N_S1_c_660_n N_A_909_74#_c_1068_n 0.0262104f $X=8.725 $Y=1.865 $X2=0
+ $Y2=0
cc_518 N_S1_c_660_n N_A_909_74#_c_1076_n 0.00102518f $X=8.725 $Y=1.865 $X2=0
+ $Y2=0
cc_519 N_S1_c_652_n N_A_909_74#_c_1071_n 8.54008e-19 $X=8.635 $Y=0.185 $X2=0
+ $Y2=0
cc_520 N_S1_M1008_g N_A_909_74#_c_1071_n 0.00120586f $X=8.71 $Y=0.92 $X2=0 $Y2=0
cc_521 N_S1_c_653_n N_VGND_c_1224_n 0.00451785f $X=7.145 $Y=0.185 $X2=0 $Y2=0
cc_522 N_S1_c_652_n N_VGND_c_1225_n 0.00308174f $X=8.635 $Y=0.185 $X2=0 $Y2=0
cc_523 N_S1_M1008_g N_VGND_c_1225_n 2.10568e-19 $X=8.71 $Y=0.92 $X2=0 $Y2=0
cc_524 N_S1_c_653_n N_VGND_c_1233_n 0.0393328f $X=7.145 $Y=0.185 $X2=0 $Y2=0
cc_525 N_S1_c_652_n N_VGND_c_1237_n 0.0409406f $X=8.635 $Y=0.185 $X2=0 $Y2=0
cc_526 N_S1_c_653_n N_VGND_c_1237_n 0.00675478f $X=7.145 $Y=0.185 $X2=0 $Y2=0
cc_527 N_A_1429_74#_c_740_n N_VPWR_M1018_d 0.00451634f $X=8.96 $Y=2.99 $X2=0
+ $Y2=0
cc_528 N_A_1429_74#_c_741_n N_VPWR_M1018_d 0.0258212f $X=9.045 $Y=2.905 $X2=0
+ $Y2=0
cc_529 N_A_1429_74#_c_740_n N_VPWR_c_836_n 0.103883f $X=8.96 $Y=2.99 $X2=0 $Y2=0
cc_530 N_A_1429_74#_c_742_n N_VPWR_c_836_n 0.0223621f $X=7.365 $Y=2.805 $X2=0
+ $Y2=0
cc_531 N_A_1429_74#_c_736_n N_VPWR_c_837_n 0.00781163f $X=9.61 $Y=1.765 $X2=0
+ $Y2=0
cc_532 N_A_1429_74#_c_730_n N_VPWR_c_837_n 0.0044907f $X=9.52 $Y=1.515 $X2=0
+ $Y2=0
cc_533 N_A_1429_74#_c_740_n N_VPWR_c_837_n 0.0142227f $X=8.96 $Y=2.99 $X2=0
+ $Y2=0
cc_534 N_A_1429_74#_c_741_n N_VPWR_c_837_n 0.0767116f $X=9.045 $Y=2.905 $X2=0
+ $Y2=0
cc_535 N_A_1429_74#_c_735_n N_VPWR_c_837_n 0.00693677f $X=9.22 $Y=1.515 $X2=0
+ $Y2=0
cc_536 N_A_1429_74#_c_737_n N_VPWR_c_839_n 0.0100916f $X=10.06 $Y=1.765 $X2=0
+ $Y2=0
cc_537 N_A_1429_74#_c_736_n N_VPWR_c_845_n 0.00422942f $X=9.61 $Y=1.765 $X2=0
+ $Y2=0
cc_538 N_A_1429_74#_c_737_n N_VPWR_c_845_n 0.00445602f $X=10.06 $Y=1.765 $X2=0
+ $Y2=0
cc_539 N_A_1429_74#_c_736_n N_VPWR_c_832_n 0.00789017f $X=9.61 $Y=1.765 $X2=0
+ $Y2=0
cc_540 N_A_1429_74#_c_737_n N_VPWR_c_832_n 0.00861067f $X=10.06 $Y=1.765 $X2=0
+ $Y2=0
cc_541 N_A_1429_74#_c_740_n N_VPWR_c_832_n 0.0597558f $X=8.96 $Y=2.99 $X2=0
+ $Y2=0
cc_542 N_A_1429_74#_c_742_n N_VPWR_c_832_n 0.0124265f $X=7.365 $Y=2.805 $X2=0
+ $Y2=0
cc_543 N_A_1429_74#_M1009_d N_A_333_74#_c_935_n 0.00411326f $X=7.145 $Y=0.37
+ $X2=0 $Y2=0
cc_544 N_A_1429_74#_c_740_n N_A_909_74#_M1017_d 0.00321405f $X=8.96 $Y=2.99
+ $X2=0 $Y2=0
cc_545 N_A_1429_74#_M1012_d N_A_909_74#_c_1072_n 0.00561204f $X=7.215 $Y=1.96
+ $X2=0 $Y2=0
cc_546 N_A_1429_74#_c_740_n N_A_909_74#_c_1072_n 0.00380094f $X=8.96 $Y=2.99
+ $X2=0 $Y2=0
cc_547 N_A_1429_74#_c_742_n N_A_909_74#_c_1072_n 0.0158897f $X=7.365 $Y=2.805
+ $X2=0 $Y2=0
cc_548 N_A_1429_74#_c_734_n N_A_909_74#_c_1066_n 0.0096883f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_549 N_A_1429_74#_M1009_d N_A_909_74#_c_1098_n 0.00481226f $X=7.145 $Y=0.37
+ $X2=0 $Y2=0
cc_550 N_A_1429_74#_c_732_n N_A_909_74#_c_1098_n 0.0134553f $X=8.96 $Y=0.34
+ $X2=0 $Y2=0
cc_551 N_A_1429_74#_c_734_n N_A_909_74#_c_1098_n 0.0198954f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_552 N_A_1429_74#_c_740_n N_A_909_74#_c_1074_n 0.0524178f $X=8.96 $Y=2.99
+ $X2=0 $Y2=0
cc_553 N_A_1429_74#_c_741_n N_A_909_74#_c_1074_n 0.0133619f $X=9.045 $Y=2.905
+ $X2=0 $Y2=0
cc_554 N_A_1429_74#_c_732_n N_A_909_74#_c_1067_n 0.0551027f $X=8.96 $Y=0.34
+ $X2=0 $Y2=0
cc_555 N_A_1429_74#_c_733_n N_A_909_74#_c_1067_n 0.00639398f $X=9.045 $Y=1.35
+ $X2=0 $Y2=0
cc_556 N_A_1429_74#_c_730_n N_A_909_74#_c_1068_n 3.30669e-19 $X=9.52 $Y=1.515
+ $X2=0 $Y2=0
cc_557 N_A_1429_74#_c_733_n N_A_909_74#_c_1068_n 0.0253617f $X=9.045 $Y=1.35
+ $X2=0 $Y2=0
cc_558 N_A_1429_74#_c_741_n N_A_909_74#_c_1068_n 0.0623724f $X=9.045 $Y=2.905
+ $X2=0 $Y2=0
cc_559 N_A_1429_74#_c_735_n N_A_909_74#_c_1068_n 0.0253857f $X=9.22 $Y=1.515
+ $X2=0 $Y2=0
cc_560 N_A_1429_74#_c_740_n N_A_909_74#_c_1076_n 0.0169546f $X=8.96 $Y=2.99
+ $X2=0 $Y2=0
cc_561 N_A_1429_74#_c_742_n N_A_909_74#_c_1076_n 0.00140699f $X=7.365 $Y=2.805
+ $X2=0 $Y2=0
cc_562 N_A_1429_74#_c_732_n N_A_909_74#_c_1071_n 0.0126013f $X=8.96 $Y=0.34
+ $X2=0 $Y2=0
cc_563 N_A_1429_74#_c_734_n N_A_909_74#_c_1071_n 2.20397e-19 $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_564 N_A_1429_74#_c_728_n X 0.0143266f $X=9.6 $Y=1.35 $X2=0 $Y2=0
cc_565 N_A_1429_74#_c_736_n X 0.00163357f $X=9.61 $Y=1.765 $X2=0 $Y2=0
cc_566 N_A_1429_74#_c_729_n X 0.0158012f $X=10.03 $Y=1.35 $X2=0 $Y2=0
cc_567 N_A_1429_74#_c_737_n X 0.00157473f $X=10.06 $Y=1.765 $X2=0 $Y2=0
cc_568 N_A_1429_74#_c_731_n X 0.0468975f $X=10.03 $Y=1.557 $X2=0 $Y2=0
cc_569 N_A_1429_74#_c_733_n X 0.00539719f $X=9.045 $Y=1.35 $X2=0 $Y2=0
cc_570 N_A_1429_74#_c_741_n X 0.00547565f $X=9.045 $Y=2.905 $X2=0 $Y2=0
cc_571 N_A_1429_74#_c_735_n X 0.0176652f $X=9.22 $Y=1.515 $X2=0 $Y2=0
cc_572 N_A_1429_74#_c_736_n X 0.00252233f $X=9.61 $Y=1.765 $X2=0 $Y2=0
cc_573 N_A_1429_74#_c_737_n X 0.00284916f $X=10.06 $Y=1.765 $X2=0 $Y2=0
cc_574 N_A_1429_74#_c_731_n X 2.74262e-19 $X=10.03 $Y=1.557 $X2=0 $Y2=0
cc_575 N_A_1429_74#_c_736_n X 0.0126237f $X=9.61 $Y=1.765 $X2=0 $Y2=0
cc_576 N_A_1429_74#_c_737_n X 0.0115887f $X=10.06 $Y=1.765 $X2=0 $Y2=0
cc_577 N_A_1429_74#_c_733_n N_VGND_M1008_d 0.0167228f $X=9.045 $Y=1.35 $X2=0
+ $Y2=0
cc_578 N_A_1429_74#_c_734_n N_VGND_c_1224_n 0.00270217f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_579 N_A_1429_74#_c_728_n N_VGND_c_1225_n 0.00403885f $X=9.6 $Y=1.35 $X2=0
+ $Y2=0
cc_580 N_A_1429_74#_c_730_n N_VGND_c_1225_n 0.00448078f $X=9.52 $Y=1.515 $X2=0
+ $Y2=0
cc_581 N_A_1429_74#_c_732_n N_VGND_c_1225_n 0.014358f $X=8.96 $Y=0.34 $X2=0
+ $Y2=0
cc_582 N_A_1429_74#_c_733_n N_VGND_c_1225_n 0.0551335f $X=9.045 $Y=1.35 $X2=0
+ $Y2=0
cc_583 N_A_1429_74#_c_735_n N_VGND_c_1225_n 0.00693677f $X=9.22 $Y=1.515 $X2=0
+ $Y2=0
cc_584 N_A_1429_74#_c_729_n N_VGND_c_1227_n 0.00577593f $X=10.03 $Y=1.35 $X2=0
+ $Y2=0
cc_585 N_A_1429_74#_c_732_n N_VGND_c_1233_n 0.105517f $X=8.96 $Y=0.34 $X2=0
+ $Y2=0
cc_586 N_A_1429_74#_c_734_n N_VGND_c_1233_n 0.0212791f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_587 N_A_1429_74#_c_728_n N_VGND_c_1234_n 0.00466874f $X=9.6 $Y=1.35 $X2=0
+ $Y2=0
cc_588 N_A_1429_74#_c_729_n N_VGND_c_1234_n 0.00466874f $X=10.03 $Y=1.35 $X2=0
+ $Y2=0
cc_589 N_A_1429_74#_c_728_n N_VGND_c_1237_n 0.00505379f $X=9.6 $Y=1.35 $X2=0
+ $Y2=0
cc_590 N_A_1429_74#_c_729_n N_VGND_c_1237_n 0.00505379f $X=10.03 $Y=1.35 $X2=0
+ $Y2=0
cc_591 N_A_1429_74#_c_732_n N_VGND_c_1237_n 0.0572698f $X=8.96 $Y=0.34 $X2=0
+ $Y2=0
cc_592 N_A_1429_74#_c_734_n N_VGND_c_1237_n 0.0110064f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_593 N_VPWR_M1004_d N_A_333_74#_c_937_n 0.00881007f $X=3.51 $Y=1.96 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_834_n N_A_333_74#_c_937_n 0.0240039f $X=3.78 $Y=2.455 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_834_n N_A_333_74#_c_972_n 0.00218589f $X=3.78 $Y=2.455 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_832_n N_A_333_74#_c_975_n 0.0261573f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_834_n N_A_333_74#_c_997_n 0.0140086f $X=3.78 $Y=2.455 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_832_n N_A_333_74#_c_997_n 0.00590416f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_599 N_VPWR_M1026_d N_A_333_74#_c_938_n 0.0103025f $X=6.18 $Y=1.96 $X2=0 $Y2=0
cc_600 N_VPWR_c_834_n N_A_333_74#_c_942_n 0.0566293f $X=3.78 $Y=2.455 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_842_n N_A_333_74#_c_942_n 0.0416012f $X=3.615 $Y=3.33 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_832_n N_A_333_74#_c_942_n 0.0338841f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_603 N_VPWR_c_844_n N_A_909_74#_c_1078_n 0.0206446f $X=6.165 $Y=3.33 $X2=0
+ $Y2=0
cc_604 N_VPWR_c_832_n N_A_909_74#_c_1078_n 0.0237181f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_605 N_VPWR_M1026_d N_A_909_74#_c_1072_n 0.00609062f $X=6.18 $Y=1.96 $X2=0
+ $Y2=0
cc_606 N_VPWR_c_835_n N_A_909_74#_c_1072_n 0.0214746f $X=6.33 $Y=2.805 $X2=0
+ $Y2=0
cc_607 N_VPWR_c_832_n N_A_909_74#_c_1072_n 0.0334778f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_608 N_VPWR_c_835_n N_A_909_74#_c_1096_n 0.0121085f $X=6.33 $Y=2.805 $X2=0
+ $Y2=0
cc_609 N_VPWR_c_844_n N_A_909_74#_c_1096_n 0.00495037f $X=6.165 $Y=3.33 $X2=0
+ $Y2=0
cc_610 N_VPWR_c_832_n N_A_909_74#_c_1096_n 0.00588467f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_611 N_VPWR_c_837_n X 0.0801844f $X=9.385 $Y=2.015 $X2=0 $Y2=0
cc_612 N_VPWR_c_839_n X 0.0781509f $X=10.285 $Y=1.985 $X2=0 $Y2=0
cc_613 N_VPWR_c_845_n X 0.0153846f $X=10.2 $Y=3.33 $X2=0 $Y2=0
cc_614 N_VPWR_c_832_n X 0.0126213f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_615 N_VPWR_c_837_n N_VGND_c_1225_n 0.00263772f $X=9.385 $Y=2.015 $X2=0 $Y2=0
cc_616 N_VPWR_c_839_n N_VGND_c_1227_n 0.00847507f $X=10.285 $Y=1.985 $X2=0 $Y2=0
cc_617 N_A_333_74#_c_937_n A_840_392# 0.00217303f $X=4.115 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_618 N_A_333_74#_c_972_n A_840_392# 0.00341048f $X=4.2 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_619 N_A_333_74#_c_975_n A_840_392# 0.0227764f $X=5.435 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_620 N_A_333_74#_c_997_n A_840_392# 6.46875e-19 $X=4.285 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_621 N_A_333_74#_c_975_n N_A_909_74#_M1015_d 0.0131238f $X=5.435 $Y=2.405
+ $X2=0 $Y2=0
cc_622 N_A_333_74#_c_939_n N_A_909_74#_M1015_d 0.00877445f $X=5.605 $Y=2.08
+ $X2=0 $Y2=0
cc_623 N_A_333_74#_c_975_n N_A_909_74#_c_1078_n 0.0233132f $X=5.435 $Y=2.405
+ $X2=0 $Y2=0
cc_624 N_A_333_74#_c_938_n N_A_909_74#_c_1078_n 0.00479616f $X=6.56 $Y=2.08
+ $X2=0 $Y2=0
cc_625 N_A_333_74#_c_939_n N_A_909_74#_c_1078_n 0.00933392f $X=5.605 $Y=2.08
+ $X2=0 $Y2=0
cc_626 N_A_333_74#_c_934_n N_A_909_74#_c_1065_n 0.010942f $X=6.73 $Y=1.195 $X2=0
+ $Y2=0
cc_627 N_A_333_74#_M1012_s N_A_909_74#_c_1072_n 0.00906302f $X=6.745 $Y=1.96
+ $X2=0 $Y2=0
cc_628 N_A_333_74#_c_938_n N_A_909_74#_c_1072_n 0.0368094f $X=6.56 $Y=2.08 $X2=0
+ $Y2=0
cc_629 N_A_333_74#_c_941_n N_A_909_74#_c_1072_n 0.021806f $X=6.9 $Y=2.115 $X2=0
+ $Y2=0
cc_630 N_A_333_74#_c_944_n N_A_909_74#_c_1072_n 0.014265f $X=6.645 $Y=2.075
+ $X2=0 $Y2=0
cc_631 N_A_333_74#_M1006_d N_A_909_74#_c_1098_n 0.00366884f $X=7.65 $Y=0.6 $X2=0
+ $Y2=0
cc_632 N_A_333_74#_c_935_n N_A_909_74#_c_1098_n 0.0520752f $X=7.79 $Y=1.195
+ $X2=0 $Y2=0
cc_633 N_A_333_74#_c_935_n N_A_909_74#_c_1073_n 0.00144295f $X=7.79 $Y=1.195
+ $X2=0 $Y2=0
cc_634 N_A_333_74#_c_941_n N_A_909_74#_c_1073_n 0.00727868f $X=6.9 $Y=2.115
+ $X2=0 $Y2=0
cc_635 N_A_333_74#_c_938_n N_A_909_74#_c_1096_n 0.0103865f $X=6.56 $Y=2.08 $X2=0
+ $Y2=0
cc_636 N_A_333_74#_c_934_n N_A_909_74#_c_1070_n 0.00365703f $X=6.73 $Y=1.195
+ $X2=0 $Y2=0
cc_637 N_A_333_74#_c_935_n N_A_909_74#_c_1070_n 0.0170427f $X=7.79 $Y=1.195
+ $X2=0 $Y2=0
cc_638 N_A_333_74#_M1006_d N_A_909_74#_c_1071_n 0.00496433f $X=7.65 $Y=0.6 $X2=0
+ $Y2=0
cc_639 N_A_333_74#_c_935_n N_A_909_74#_c_1071_n 0.00845717f $X=7.79 $Y=1.195
+ $X2=0 $Y2=0
cc_640 N_A_333_74#_c_938_n A_1152_392# 0.00623161f $X=6.56 $Y=2.08 $X2=-0.19
+ $Y2=-0.245
cc_641 N_A_333_74#_c_946_n A_507_74# 0.00418009f $X=2.495 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_642 N_A_909_74#_c_1072_n A_1152_392# 0.0012425f $X=7.65 $Y=2.455 $X2=-0.19
+ $Y2=-0.245
cc_643 N_A_909_74#_c_1096_n A_1152_392# 0.00742261f $X=5.86 $Y=2.455 $X2=-0.19
+ $Y2=-0.245
cc_644 N_A_909_74#_c_1065_n N_VGND_M1011_d 0.00832719f $X=6.69 $Y=0.855 $X2=0
+ $Y2=0
cc_645 N_A_909_74#_c_1069_n N_VGND_c_1223_n 0.01805f $X=4.855 $Y=0.515 $X2=0
+ $Y2=0
cc_646 N_A_909_74#_c_1065_n N_VGND_c_1224_n 0.0213424f $X=6.69 $Y=0.855 $X2=0
+ $Y2=0
cc_647 N_A_909_74#_c_1066_n N_VGND_c_1224_n 0.0170237f $X=6.855 $Y=0.515 $X2=0
+ $Y2=0
cc_648 N_A_909_74#_c_1069_n N_VGND_c_1230_n 0.0252084f $X=4.855 $Y=0.515 $X2=0
+ $Y2=0
cc_649 N_A_909_74#_c_1066_n N_VGND_c_1233_n 0.0109523f $X=6.855 $Y=0.515 $X2=0
+ $Y2=0
cc_650 N_A_909_74#_c_1065_n N_VGND_c_1237_n 0.0454954f $X=6.69 $Y=0.855 $X2=0
+ $Y2=0
cc_651 N_A_909_74#_c_1066_n N_VGND_c_1237_n 0.00911557f $X=6.855 $Y=0.515 $X2=0
+ $Y2=0
cc_652 N_A_909_74#_c_1098_n N_VGND_c_1237_n 0.00732805f $X=7.845 $Y=0.855 $X2=0
+ $Y2=0
cc_653 N_A_909_74#_c_1069_n N_VGND_c_1237_n 0.0209023f $X=4.855 $Y=0.515 $X2=0
+ $Y2=0
cc_654 N_A_909_74#_c_1065_n A_1047_74# 0.0266143f $X=6.69 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_655 X N_VGND_c_1225_n 0.0286545f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_656 X N_VGND_c_1227_n 0.0323784f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_657 X N_VGND_c_1234_n 0.0105983f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_658 X N_VGND_c_1237_n 0.0113894f $X=9.755 $Y=0.47 $X2=0 $Y2=0
