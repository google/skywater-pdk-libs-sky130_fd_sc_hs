* File: sky130_fd_sc_hs__or4b_1.pxi.spice
* Created: Tue Sep  1 20:21:22 2020
* 
x_PM_SKY130_FD_SC_HS__OR4B_1%D_N N_D_N_M1008_g N_D_N_c_81_n N_D_N_c_84_n
+ N_D_N_c_85_n N_D_N_M1004_g D_N N_D_N_c_82_n PM_SKY130_FD_SC_HS__OR4B_1%D_N
x_PM_SKY130_FD_SC_HS__OR4B_1%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1004_s
+ N_A_27_74#_M1010_g N_A_27_74#_c_118_n N_A_27_74#_c_126_n N_A_27_74#_M1009_g
+ N_A_27_74#_c_119_n N_A_27_74#_c_127_n N_A_27_74#_c_120_n N_A_27_74#_c_121_n
+ N_A_27_74#_c_128_n N_A_27_74#_c_129_n N_A_27_74#_c_122_n N_A_27_74#_c_123_n
+ N_A_27_74#_c_124_n PM_SKY130_FD_SC_HS__OR4B_1%A_27_74#
x_PM_SKY130_FD_SC_HS__OR4B_1%C N_C_c_189_n N_C_c_194_n N_C_M1005_g N_C_M1002_g C
+ C N_C_c_190_n N_C_c_191_n N_C_c_192_n PM_SKY130_FD_SC_HS__OR4B_1%C
x_PM_SKY130_FD_SC_HS__OR4B_1%B N_B_c_226_n N_B_c_231_n N_B_M1007_g N_B_M1006_g B
+ B N_B_c_229_n PM_SKY130_FD_SC_HS__OR4B_1%B
x_PM_SKY130_FD_SC_HS__OR4B_1%A N_A_c_262_n N_A_M1000_g N_A_M1011_g A N_A_c_264_n
+ PM_SKY130_FD_SC_HS__OR4B_1%A
x_PM_SKY130_FD_SC_HS__OR4B_1%A_228_74# N_A_228_74#_M1010_d N_A_228_74#_M1006_d
+ N_A_228_74#_M1009_s N_A_228_74#_c_301_n N_A_228_74#_M1001_g
+ N_A_228_74#_M1003_g N_A_228_74#_c_313_n N_A_228_74#_c_303_n
+ N_A_228_74#_c_310_n N_A_228_74#_c_331_n N_A_228_74#_c_322_n
+ N_A_228_74#_c_304_n N_A_228_74#_c_305_n N_A_228_74#_c_306_n
+ N_A_228_74#_c_307_n N_A_228_74#_c_312_n PM_SKY130_FD_SC_HS__OR4B_1%A_228_74#
x_PM_SKY130_FD_SC_HS__OR4B_1%VPWR N_VPWR_M1004_d N_VPWR_M1000_d N_VPWR_c_402_n
+ N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n VPWR N_VPWR_c_406_n
+ N_VPWR_c_407_n N_VPWR_c_401_n N_VPWR_c_409_n PM_SKY130_FD_SC_HS__OR4B_1%VPWR
x_PM_SKY130_FD_SC_HS__OR4B_1%X N_X_M1003_d N_X_M1001_d N_X_c_445_n N_X_c_446_n X
+ X X X N_X_c_447_n PM_SKY130_FD_SC_HS__OR4B_1%X
x_PM_SKY130_FD_SC_HS__OR4B_1%VGND N_VGND_M1008_d N_VGND_M1002_d N_VGND_M1011_d
+ N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n
+ N_VGND_c_476_n N_VGND_c_477_n VGND N_VGND_c_478_n N_VGND_c_479_n
+ N_VGND_c_480_n N_VGND_c_481_n PM_SKY130_FD_SC_HS__OR4B_1%VGND
cc_1 VNB N_D_N_M1008_g 0.0540783f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_D_N_c_81_n 0.0220576f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.78
cc_3 VNB N_D_N_c_82_n 0.0105114f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_4 VNB N_A_27_74#_M1010_g 0.0569092f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_5 VNB N_A_27_74#_c_118_n 0.029762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_74#_c_119_n 0.0322397f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_7 VNB N_A_27_74#_c_120_n 0.0122485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_121_n 0.0101326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_122_n 0.00550808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_123_n 0.00125837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_124_n 0.0097753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_c_189_n 0.01609f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_13 VNB N_C_c_190_n 0.0339822f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_14 VNB N_C_c_191_n 0.0111854f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_15 VNB N_C_c_192_n 0.0244906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_226_n 0.00788532f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_17 VNB N_B_M1006_g 0.0275918f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_18 VNB B 0.0044004f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_B_c_229_n 0.0327832f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_20 VNB N_A_c_262_n 0.0275752f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_21 VNB N_A_M1011_g 0.0361617f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.955
cc_22 VNB N_A_c_264_n 0.00165719f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.615
cc_23 VNB N_A_228_74#_c_301_n 0.0363572f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_228_74#_M1003_g 0.0294785f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_25 VNB N_A_228_74#_c_303_n 0.0177655f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_26 VNB N_A_228_74#_c_304_n 0.0139115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_228_74#_c_305_n 0.0110547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_228_74#_c_306_n 0.0112948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_228_74#_c_307_n 3.99197e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_401_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_445_n 0.0272846f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_32 VNB N_X_c_446_n 0.0154926f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_33 VNB N_X_c_447_n 0.0248107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_471_n 0.01314f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.615
cc_35 VNB N_VGND_c_472_n 0.00984011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_473_n 0.00981014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_474_n 0.0365984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_475_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_476_n 0.0195351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_477_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_478_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_479_n 0.0211504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_480_n 0.258711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_481_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_D_N_c_81_n 0.0143306f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.78
cc_46 VPB N_D_N_c_84_n 0.0144478f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.955
cc_47 VPB N_D_N_c_85_n 0.0287331f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.045
cc_48 VPB N_D_N_c_82_n 0.00566928f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_49 VPB N_A_27_74#_c_118_n 0.0267234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_27_74#_c_126_n 0.0167678f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_51 VPB N_A_27_74#_c_127_n 0.0353617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_27_74#_c_128_n 0.00616913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_74#_c_129_n 0.00989919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_74#_c_123_n 0.0133601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_74#_c_124_n 0.0236232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_C_c_189_n 5.92781e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_57 VPB N_C_c_194_n 0.0196169f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_58 VPB N_C_c_191_n 0.00377678f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_59 VPB N_B_c_226_n 7.40903e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_60 VPB N_B_c_231_n 0.0214257f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_61 VPB B 0.00255974f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_62 VPB N_A_c_262_n 0.0293416f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_63 VPB N_A_c_264_n 0.00244101f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.615
cc_64 VPB N_A_228_74#_c_301_n 0.0299331f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_65 VPB N_A_228_74#_c_303_n 0.00136231f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_66 VPB N_A_228_74#_c_310_n 0.0173855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_228_74#_c_307_n 0.00301535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_228_74#_c_312_n 0.00218793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_402_n 0.0211975f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.54
cc_70 VPB N_VPWR_c_403_n 0.0143486f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_71 VPB N_VPWR_c_404_n 0.0738078f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_72 VPB N_VPWR_c_405_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_406_n 0.0192906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_407_n 0.0198775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_401_n 0.127348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_409_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB X 0.0155822f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_78 VPB X 0.0431281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_X_c_447_n 0.00761759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 N_D_N_M1008_g N_A_27_74#_M1010_g 0.0285007f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_81 N_D_N_M1008_g N_A_27_74#_c_119_n 0.017246f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_82 N_D_N_c_85_n N_A_27_74#_c_127_n 0.0178576f $X=0.51 $Y=2.045 $X2=0 $Y2=0
cc_83 N_D_N_M1008_g N_A_27_74#_c_120_n 0.0115704f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_84 N_D_N_c_81_n N_A_27_74#_c_120_n 7.18829e-19 $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_85 N_D_N_c_82_n N_A_27_74#_c_120_n 0.00889268f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_86 N_D_N_M1008_g N_A_27_74#_c_121_n 0.00419718f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_87 N_D_N_c_81_n N_A_27_74#_c_121_n 0.00419322f $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_88 N_D_N_c_82_n N_A_27_74#_c_121_n 0.0273487f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_89 N_D_N_c_84_n N_A_27_74#_c_128_n 0.00238554f $X=0.51 $Y=1.955 $X2=0 $Y2=0
cc_90 N_D_N_c_85_n N_A_27_74#_c_128_n 0.0118217f $X=0.51 $Y=2.045 $X2=0 $Y2=0
cc_91 N_D_N_c_82_n N_A_27_74#_c_128_n 0.00853562f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_92 N_D_N_c_81_n N_A_27_74#_c_129_n 0.00419322f $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_93 N_D_N_c_84_n N_A_27_74#_c_129_n 4.3488e-19 $X=0.51 $Y=1.955 $X2=0 $Y2=0
cc_94 N_D_N_c_85_n N_A_27_74#_c_129_n 0.00403309f $X=0.51 $Y=2.045 $X2=0 $Y2=0
cc_95 N_D_N_c_82_n N_A_27_74#_c_129_n 0.0277478f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_96 N_D_N_M1008_g N_A_27_74#_c_122_n 0.00344365f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_97 N_D_N_c_81_n N_A_27_74#_c_122_n 4.69863e-19 $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_98 N_D_N_c_82_n N_A_27_74#_c_122_n 0.00765956f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_99 N_D_N_c_81_n N_A_27_74#_c_123_n 0.00149088f $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_100 N_D_N_c_84_n N_A_27_74#_c_123_n 0.00134246f $X=0.51 $Y=1.955 $X2=0 $Y2=0
cc_101 N_D_N_c_82_n N_A_27_74#_c_123_n 0.0116895f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_102 N_D_N_c_81_n N_A_27_74#_c_124_n 0.0200876f $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_103 N_D_N_c_82_n N_A_27_74#_c_124_n 2.41258e-19 $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_104 N_D_N_c_85_n N_VPWR_c_402_n 0.018269f $X=0.51 $Y=2.045 $X2=0 $Y2=0
cc_105 N_D_N_c_85_n N_VPWR_c_406_n 0.00445602f $X=0.51 $Y=2.045 $X2=0 $Y2=0
cc_106 N_D_N_c_85_n N_VPWR_c_401_n 0.0086523f $X=0.51 $Y=2.045 $X2=0 $Y2=0
cc_107 N_D_N_M1008_g N_VGND_c_471_n 0.00689618f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_108 N_D_N_M1008_g N_VGND_c_478_n 0.00434272f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_109 N_D_N_M1008_g N_VGND_c_480_n 0.0082497f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_110 N_A_27_74#_c_118_n N_C_c_189_n 0.00822497f $X=1.63 $Y=1.69 $X2=0 $Y2=0
cc_111 N_A_27_74#_c_126_n N_C_c_194_n 0.0575646f $X=1.705 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_27_74#_c_118_n N_C_c_191_n 0.00137289f $X=1.63 $Y=1.69 $X2=0 $Y2=0
cc_113 N_A_27_74#_M1010_g N_A_228_74#_c_313_n 0.00500409f $X=1.065 $Y=0.645
+ $X2=0 $Y2=0
cc_114 N_A_27_74#_M1010_g N_A_228_74#_c_303_n 0.0172544f $X=1.065 $Y=0.645 $X2=0
+ $Y2=0
cc_115 N_A_27_74#_c_118_n N_A_228_74#_c_303_n 0.023702f $X=1.63 $Y=1.69 $X2=0
+ $Y2=0
cc_116 N_A_27_74#_c_126_n N_A_228_74#_c_303_n 0.00416376f $X=1.705 $Y=1.765
+ $X2=0 $Y2=0
cc_117 N_A_27_74#_c_120_n N_A_228_74#_c_303_n 0.00935581f $X=0.81 $Y=1.195 $X2=0
+ $Y2=0
cc_118 N_A_27_74#_c_122_n N_A_228_74#_c_303_n 0.0147829f $X=0.895 $Y=1.58 $X2=0
+ $Y2=0
cc_119 N_A_27_74#_c_123_n N_A_228_74#_c_303_n 0.0270211f $X=0.975 $Y=1.745 $X2=0
+ $Y2=0
cc_120 N_A_27_74#_c_124_n N_A_228_74#_c_303_n 8.53863e-19 $X=0.975 $Y=1.69 $X2=0
+ $Y2=0
cc_121 N_A_27_74#_c_126_n N_A_228_74#_c_310_n 0.0134092f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_27_74#_c_126_n N_A_228_74#_c_322_n 0.015358f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_27_74#_c_126_n N_A_228_74#_c_312_n 2.24111e-19 $X=1.705 $Y=1.765
+ $X2=0 $Y2=0
cc_124 N_A_27_74#_c_123_n N_A_228_74#_c_312_n 0.00991941f $X=0.975 $Y=1.745
+ $X2=0 $Y2=0
cc_125 N_A_27_74#_c_123_n N_VPWR_M1004_d 0.00132795f $X=0.975 $Y=1.745 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_27_74#_c_126_n N_VPWR_c_402_n 0.00364201f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A_27_74#_c_127_n N_VPWR_c_402_n 0.0266809f $X=0.285 $Y=2.265 $X2=0
+ $Y2=0
cc_128 N_A_27_74#_c_128_n N_VPWR_c_402_n 0.014648f $X=0.81 $Y=2.035 $X2=0 $Y2=0
cc_129 N_A_27_74#_c_123_n N_VPWR_c_402_n 0.0125996f $X=0.975 $Y=1.745 $X2=0
+ $Y2=0
cc_130 N_A_27_74#_c_124_n N_VPWR_c_402_n 6.80259e-19 $X=0.975 $Y=1.69 $X2=0
+ $Y2=0
cc_131 N_A_27_74#_c_126_n N_VPWR_c_404_n 0.00481995f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_27_74#_c_127_n N_VPWR_c_406_n 0.0145938f $X=0.285 $Y=2.265 $X2=0
+ $Y2=0
cc_133 N_A_27_74#_c_126_n N_VPWR_c_401_n 0.00508379f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A_27_74#_c_127_n N_VPWR_c_401_n 0.0120466f $X=0.285 $Y=2.265 $X2=0
+ $Y2=0
cc_135 N_A_27_74#_M1010_g N_VGND_c_471_n 0.00733509f $X=1.065 $Y=0.645 $X2=0
+ $Y2=0
cc_136 N_A_27_74#_c_119_n N_VGND_c_471_n 0.0237192f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_137 N_A_27_74#_c_120_n N_VGND_c_471_n 0.028903f $X=0.81 $Y=1.195 $X2=0 $Y2=0
cc_138 N_A_27_74#_c_124_n N_VGND_c_471_n 4.14455e-19 $X=0.975 $Y=1.69 $X2=0
+ $Y2=0
cc_139 N_A_27_74#_M1010_g N_VGND_c_474_n 0.00437222f $X=1.065 $Y=0.645 $X2=0
+ $Y2=0
cc_140 N_A_27_74#_c_119_n N_VGND_c_478_n 0.0145639f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_141 N_A_27_74#_M1010_g N_VGND_c_480_n 0.00828236f $X=1.065 $Y=0.645 $X2=0
+ $Y2=0
cc_142 N_A_27_74#_c_119_n N_VGND_c_480_n 0.0119984f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_143 N_C_c_189_n N_B_c_226_n 0.0100481f $X=2.125 $Y=1.675 $X2=0 $Y2=0
cc_144 N_C_c_194_n N_B_c_231_n 0.0722811f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_145 N_C_c_191_n N_B_M1006_g 0.00276524f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_146 N_C_c_192_n N_B_M1006_g 0.0209778f $X=2.05 $Y=1.045 $X2=0 $Y2=0
cc_147 N_C_c_190_n B 6.63977e-19 $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_148 N_C_c_191_n B 0.0460922f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_149 N_C_c_190_n N_B_c_229_n 0.0100481f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_150 N_C_c_191_n N_B_c_229_n 0.00348274f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_151 N_C_c_189_n N_A_228_74#_c_303_n 0.00135712f $X=2.125 $Y=1.675 $X2=0 $Y2=0
cc_152 N_C_c_194_n N_A_228_74#_c_303_n 8.25834e-19 $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_153 N_C_c_190_n N_A_228_74#_c_303_n 0.00720024f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_154 N_C_c_191_n N_A_228_74#_c_303_n 0.0465537f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_155 N_C_c_192_n N_A_228_74#_c_303_n 0.00442451f $X=2.05 $Y=1.045 $X2=0 $Y2=0
cc_156 N_C_c_194_n N_A_228_74#_c_310_n 0.00355341f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_157 N_C_c_190_n N_A_228_74#_c_331_n 0.00117855f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_158 N_C_c_191_n N_A_228_74#_c_331_n 0.0144123f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_159 N_C_c_192_n N_A_228_74#_c_331_n 0.00417451f $X=2.05 $Y=1.045 $X2=0 $Y2=0
cc_160 N_C_c_194_n N_A_228_74#_c_322_n 0.0148544f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_161 N_C_c_190_n N_A_228_74#_c_322_n 4.10942e-19 $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_162 N_C_c_191_n N_A_228_74#_c_322_n 0.0270527f $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_163 N_C_c_192_n N_A_228_74#_c_304_n 3.19871e-19 $X=2.05 $Y=1.045 $X2=0 $Y2=0
cc_164 N_C_c_194_n N_VPWR_c_404_n 0.0049405f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_165 N_C_c_194_n N_VPWR_c_401_n 0.00508379f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_166 N_C_c_191_n N_VGND_c_472_n 6.99196e-19 $X=2.05 $Y=1.21 $X2=0 $Y2=0
cc_167 N_C_c_192_n N_VGND_c_472_n 0.00681565f $X=2.05 $Y=1.045 $X2=0 $Y2=0
cc_168 N_C_c_192_n N_VGND_c_474_n 0.00437241f $X=2.05 $Y=1.045 $X2=0 $Y2=0
cc_169 N_C_c_192_n N_VGND_c_480_n 0.00828273f $X=2.05 $Y=1.045 $X2=0 $Y2=0
cc_170 N_B_c_226_n N_A_c_262_n 0.00765573f $X=2.545 $Y=1.675 $X2=-0.19
+ $Y2=-0.245
cc_171 N_B_c_231_n N_A_c_262_n 0.043694f $X=2.545 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_172 B N_A_c_262_n 0.00247286f $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_173 N_B_c_229_n N_A_c_262_n 0.0097505f $X=2.62 $Y=1.345 $X2=-0.19 $Y2=-0.245
cc_174 N_B_M1006_g N_A_M1011_g 0.0314674f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_175 B N_A_M1011_g 0.00106272f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_176 N_B_c_226_n N_A_c_264_n 2.61717e-19 $X=2.545 $Y=1.675 $X2=0 $Y2=0
cc_177 B N_A_c_264_n 0.0284474f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_178 N_B_c_229_n N_A_c_264_n 5.57265e-19 $X=2.62 $Y=1.345 $X2=0 $Y2=0
cc_179 N_B_c_231_n N_A_228_74#_c_322_n 0.015481f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_180 B N_A_228_74#_c_322_n 0.0233594f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_181 N_B_c_229_n N_A_228_74#_c_322_n 5.11979e-19 $X=2.62 $Y=1.345 $X2=0 $Y2=0
cc_182 N_B_M1006_g N_A_228_74#_c_304_n 0.0158484f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_183 B N_A_228_74#_c_304_n 0.00150773f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_184 N_B_c_231_n N_VPWR_c_404_n 0.0049405f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_185 N_B_c_231_n N_VPWR_c_401_n 0.00508379f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_186 N_B_M1006_g N_VGND_c_472_n 0.00643859f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_187 B N_VGND_c_472_n 0.00700995f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_188 N_B_c_229_n N_VGND_c_472_n 9.27026e-19 $X=2.62 $Y=1.345 $X2=0 $Y2=0
cc_189 N_B_M1006_g N_VGND_c_476_n 0.00434272f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_190 N_B_M1006_g N_VGND_c_480_n 0.0082141f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_191 N_A_c_262_n N_A_228_74#_c_301_n 0.0352503f $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_M1011_g N_A_228_74#_c_301_n 0.00152487f $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_193 N_A_c_264_n N_A_228_74#_c_301_n 3.09225e-19 $X=3.16 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A_M1011_g N_A_228_74#_M1003_g 0.0170961f $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_195 N_A_c_262_n N_A_228_74#_c_322_n 0.0172667f $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_c_264_n N_A_228_74#_c_322_n 0.0226548f $X=3.16 $Y=1.515 $X2=0 $Y2=0
cc_197 N_A_c_262_n N_A_228_74#_c_304_n 5.40529e-19 $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A_M1011_g N_A_228_74#_c_304_n 0.0165678f $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_199 N_A_c_264_n N_A_228_74#_c_304_n 0.0108629f $X=3.16 $Y=1.515 $X2=0 $Y2=0
cc_200 N_A_c_262_n N_A_228_74#_c_305_n 7.68393e-19 $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_M1011_g N_A_228_74#_c_305_n 0.00931685f $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_202 N_A_c_264_n N_A_228_74#_c_305_n 0.0149678f $X=3.16 $Y=1.515 $X2=0 $Y2=0
cc_203 N_A_c_262_n N_A_228_74#_c_306_n 0.00172222f $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A_M1011_g N_A_228_74#_c_306_n 0.00349438f $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_205 N_A_c_264_n N_A_228_74#_c_306_n 0.022612f $X=3.16 $Y=1.515 $X2=0 $Y2=0
cc_206 N_A_c_262_n N_A_228_74#_c_307_n 0.00381314f $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A_c_264_n N_A_228_74#_c_307_n 0.0116479f $X=3.16 $Y=1.515 $X2=0 $Y2=0
cc_208 N_A_c_262_n N_VPWR_c_403_n 0.0176002f $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A_c_262_n N_VPWR_c_404_n 0.0049405f $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_c_262_n N_VPWR_c_401_n 0.00508379f $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A_M1011_g N_X_c_445_n 8.4339e-19 $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_212 N_A_c_262_n X 8.15898e-19 $X=3.085 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A_M1011_g N_VGND_c_473_n 0.00780925f $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_214 N_A_M1011_g N_VGND_c_476_n 0.00394617f $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_215 N_A_M1011_g N_VGND_c_480_n 0.00694298f $X=3.14 $Y=0.645 $X2=0 $Y2=0
cc_216 N_A_228_74#_c_322_n N_VPWR_M1000_d 0.0180857f $X=3.495 $Y=2.035 $X2=0
+ $Y2=0
cc_217 N_A_228_74#_c_307_n N_VPWR_M1000_d 0.00232437f $X=3.58 $Y=1.95 $X2=0
+ $Y2=0
cc_218 N_A_228_74#_c_310_n N_VPWR_c_402_n 0.0279895f $X=1.48 $Y=2.695 $X2=0
+ $Y2=0
cc_219 N_A_228_74#_c_301_n N_VPWR_c_403_n 0.0103777f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_220 N_A_228_74#_c_322_n N_VPWR_c_403_n 0.0261984f $X=3.495 $Y=2.035 $X2=0
+ $Y2=0
cc_221 N_A_228_74#_c_310_n N_VPWR_c_404_n 0.0097982f $X=1.48 $Y=2.695 $X2=0
+ $Y2=0
cc_222 N_A_228_74#_c_301_n N_VPWR_c_407_n 0.00445602f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_A_228_74#_c_301_n N_VPWR_c_401_n 0.00865339f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_224 N_A_228_74#_c_310_n N_VPWR_c_401_n 0.0111907f $X=1.48 $Y=2.695 $X2=0
+ $Y2=0
cc_225 N_A_228_74#_c_322_n A_356_368# 0.00885531f $X=3.495 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_228_74#_c_322_n A_440_368# 0.0114366f $X=3.495 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_228_74#_c_322_n A_524_368# 0.0182491f $X=3.495 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_228_74#_M1003_g N_X_c_445_n 0.0094414f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A_228_74#_c_301_n N_X_c_446_n 2.76807e-19 $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A_228_74#_M1003_g N_X_c_446_n 0.00374195f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_228_74#_c_306_n N_X_c_446_n 0.0104426f $X=3.58 $Y=1.63 $X2=0 $Y2=0
cc_232 N_A_228_74#_c_301_n X 0.00325705f $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_228_74#_c_306_n X 0.00453218f $X=3.58 $Y=1.63 $X2=0 $Y2=0
cc_234 N_A_228_74#_c_307_n X 0.00573847f $X=3.58 $Y=1.95 $X2=0 $Y2=0
cc_235 N_A_228_74#_c_301_n X 0.0130205f $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A_228_74#_c_301_n N_X_c_447_n 0.005314f $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_228_74#_M1003_g N_X_c_447_n 0.00246301f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_228_74#_c_306_n N_X_c_447_n 0.0302873f $X=3.58 $Y=1.63 $X2=0 $Y2=0
cc_239 N_A_228_74#_c_307_n N_X_c_447_n 0.00578887f $X=3.58 $Y=1.95 $X2=0 $Y2=0
cc_240 N_A_228_74#_c_305_n N_VGND_M1011_d 5.47736e-19 $X=3.495 $Y=1.095 $X2=0
+ $Y2=0
cc_241 N_A_228_74#_c_306_n N_VGND_M1011_d 0.00361029f $X=3.58 $Y=1.63 $X2=0
+ $Y2=0
cc_242 N_A_228_74#_c_303_n N_VGND_c_471_n 0.00193998f $X=1.48 $Y=1.95 $X2=0
+ $Y2=0
cc_243 N_A_228_74#_c_304_n N_VGND_c_472_n 0.0162996f $X=2.942 $Y=0.758 $X2=0
+ $Y2=0
cc_244 N_A_228_74#_c_301_n N_VGND_c_473_n 2.48813e-19 $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_245 N_A_228_74#_M1003_g N_VGND_c_473_n 0.00805958f $X=3.785 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_228_74#_c_304_n N_VGND_c_473_n 0.0383459f $X=2.942 $Y=0.758 $X2=0
+ $Y2=0
cc_247 N_A_228_74#_c_305_n N_VGND_c_473_n 0.0163722f $X=3.495 $Y=1.095 $X2=0
+ $Y2=0
cc_248 N_A_228_74#_c_306_n N_VGND_c_473_n 0.0116309f $X=3.58 $Y=1.63 $X2=0 $Y2=0
cc_249 N_A_228_74#_c_313_n N_VGND_c_474_n 0.0117263f $X=1.48 $Y=0.875 $X2=0
+ $Y2=0
cc_250 N_A_228_74#_c_331_n N_VGND_c_474_n 0.00939361f $X=1.925 $Y=0.71 $X2=0
+ $Y2=0
cc_251 N_A_228_74#_c_304_n N_VGND_c_476_n 0.0158618f $X=2.942 $Y=0.758 $X2=0
+ $Y2=0
cc_252 N_A_228_74#_M1003_g N_VGND_c_479_n 0.00434272f $X=3.785 $Y=0.74 $X2=0
+ $Y2=0
cc_253 N_A_228_74#_M1003_g N_VGND_c_480_n 0.00826503f $X=3.785 $Y=0.74 $X2=0
+ $Y2=0
cc_254 N_A_228_74#_c_313_n N_VGND_c_480_n 0.0168429f $X=1.48 $Y=0.875 $X2=0
+ $Y2=0
cc_255 N_A_228_74#_c_331_n N_VGND_c_480_n 0.0138323f $X=1.925 $Y=0.71 $X2=0
+ $Y2=0
cc_256 N_A_228_74#_c_304_n N_VGND_c_480_n 0.0129722f $X=2.942 $Y=0.758 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_403_n X 0.0274544f $X=3.5 $Y=2.455 $X2=0 $Y2=0
cc_258 N_VPWR_c_407_n X 0.0177173f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_259 N_VPWR_c_401_n X 0.0146319f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_260 N_X_c_445_n N_VGND_c_473_n 0.0328261f $X=4 $Y=0.515 $X2=0 $Y2=0
cc_261 N_X_c_445_n N_VGND_c_479_n 0.0176874f $X=4 $Y=0.515 $X2=0 $Y2=0
cc_262 N_X_c_445_n N_VGND_c_480_n 0.0145837f $X=4 $Y=0.515 $X2=0 $Y2=0
