* File: sky130_fd_sc_hs__dfrtp_1.pex.spice
* Created: Tue Sep  1 19:59:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFRTP_1%D 2 4 5 7 10 12 13 14 19 20 23
r32 23 25 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.845
+ $X2=0.402 $Y2=2.01
r33 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r34 19 21 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.165
+ $X2=0.402 $Y2=1
r35 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r36 14 24 5.61447 $w=3.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.32 $Y=2.035
+ $X2=0.32 $Y2=1.845
r37 13 24 5.31897 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.32 $Y=1.665
+ $X2=0.32 $Y2=1.845
r38 12 13 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.665
r39 12 20 3.84148 $w=3.88e-07 $l=1.3e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.165
r40 10 21 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.51 $Y=0.6 $X2=0.51
+ $Y2=1
r41 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=2.465
+ $X2=0.495 $Y2=2.75
r42 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=2.375 $X2=0.495
+ $Y2=2.465
r43 4 25 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=0.495 $Y=2.375
+ $X2=0.495 $Y2=2.01
r44 2 23 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.828
+ $X2=0.402 $Y2=1.845
r45 1 19 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.165
r46 1 2 102.129 $w=3.65e-07 $l=6.46e-07 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.828
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%RESET_B 3 6 8 9 11 12 14 15 17 19 22 24 26
+ 29 31 32 33 34 37 39 42 45 46 49 53 59
c201 46 0 1.47238e-19 $X=1.155 $Y=1.295
c202 45 0 1.09291e-19 $X=1.155 $Y=1.295
c203 33 0 3.91908e-20 $X=7.775 $Y=2.035
c204 29 0 9.2224e-20 $X=4.875 $Y=1.26
c205 12 0 1.54159e-19 $X=4.785 $Y=1.185
r206 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.18
+ $Y=2.09 $X2=8.18 $Y2=2.09
r207 53 55 32.8941 $w=3.59e-07 $l=2.45e-07 $layer=POLY_cond $X=4.875 $Y=2.002
+ $X2=5.12 $Y2=2.002
r208 52 53 2.01393 $w=3.59e-07 $l=1.5e-08 $layer=POLY_cond $X=4.86 $Y=2.002
+ $X2=4.875 $Y2=2.002
r209 49 51 40.6549 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.072 $Y=1.975
+ $X2=1.072 $Y2=2.14
r210 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.975 $X2=1.155 $Y2=1.975
r211 46 50 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.975
r212 45 47 46.3954 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.072 $Y=1.295
+ $X2=1.072 $Y2=1.13
r213 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.295 $X2=1.155 $Y2=1.295
r214 42 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r215 40 59 8.94433 $w=3.33e-07 $l=2.6e-07 $layer=LI1_cond $X=7.92 $Y=2.087
+ $X2=8.18 $Y2=2.087
r216 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r217 37 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.96 $X2=5.12 $Y2=1.96
r218 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r219 34 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=2.035
+ $X2=5.04 $Y2=2.035
r220 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r221 33 34 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.185 $Y2=2.035
r222 32 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r223 31 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r224 31 32 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=1.345 $Y2=2.035
r225 27 29 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.785 $Y=1.26
+ $X2=4.875 $Y2=1.26
r226 24 58 61.0536 $w=2.9e-07 $l=3.36749e-07 $layer=POLY_cond $X=8.26 $Y=2.39
+ $X2=8.182 $Y2=2.09
r227 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.26 $Y=2.39
+ $X2=8.26 $Y2=2.675
r228 20 58 38.6157 $w=2.9e-07 $l=1.76125e-07 $layer=POLY_cond $X=8.205 $Y=1.925
+ $X2=8.182 $Y2=2.09
r229 20 22 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=8.205 $Y=1.925
+ $X2=8.205 $Y2=0.615
r230 19 53 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.875 $Y=1.795
+ $X2=4.875 $Y2=2.002
r231 18 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.875 $Y=1.335
+ $X2=4.875 $Y2=1.26
r232 18 19 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.875 $Y=1.335
+ $X2=4.875 $Y2=1.795
r233 15 52 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.86 $Y=2.21
+ $X2=4.86 $Y2=2.002
r234 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.86 $Y=2.21
+ $X2=4.86 $Y2=2.495
r235 12 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.785 $Y=1.185
+ $X2=4.785 $Y2=1.26
r236 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.785 $Y=1.185
+ $X2=4.785 $Y2=0.9
r237 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.945 $Y=2.465
+ $X2=0.945 $Y2=2.75
r238 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.945 $Y=2.375
+ $X2=0.945 $Y2=2.465
r239 8 51 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.945 $Y=2.375
+ $X2=0.945 $Y2=2.14
r240 6 49 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=1.072 $Y=1.893
+ $X2=1.072 $Y2=1.975
r241 5 45 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=1.072 $Y=1.377
+ $X2=1.072 $Y2=1.295
r242 5 6 55.7728 $w=4.95e-07 $l=5.16e-07 $layer=POLY_cond $X=1.072 $Y=1.377
+ $X2=1.072 $Y2=1.893
r243 3 47 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.9 $Y=0.6 $X2=0.9
+ $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%CLK 3 5 7 8
c43 5 0 3.04755e-19 $X=1.925 $Y=1.755
c44 3 0 7.58493e-21 $X=1.89 $Y=0.74
r45 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.475 $X2=1.91 $Y2=1.475
r46 8 12 7.68262 $w=3.97e-07 $l=2.5e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.91 $Y2=1.545
r47 5 11 57.6553 $w=2.91e-07 $l=2.87402e-07 $layer=POLY_cond $X=1.925 $Y=1.755
+ $X2=1.91 $Y2=1.475
r48 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.925 $Y=1.755
+ $X2=1.925 $Y2=2.39
r49 1 11 38.6072 $w=2.91e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.89 $Y=1.31
+ $X2=1.91 $Y2=1.475
r50 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.89 $Y=1.31 $X2=1.89
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%A_490_366# 1 2 8 9 11 12 14 16 18 20 21 22
+ 23 25 29 32 33 35 37 40 43 44 45 48 52 53 60 66 69 71
c201 60 0 1.33783e-19 $X=4.35 $Y=0.415
c202 43 0 2.03762e-20 $X=5.565 $Y=0.565
c203 22 0 1.83796e-19 $X=6.33 $Y=1.27
c204 16 0 1.00917e-19 $X=4.005 $Y=0.9
r205 68 69 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=7.13 $Y=1.18
+ $X2=7.335 $Y2=1.18
r206 66 77 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.855 $Y=1.18
+ $X2=6.855 $Y2=1.27
r207 65 68 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.855 $Y=1.18
+ $X2=7.13 $Y2=1.18
r208 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.855
+ $Y=1.18 $X2=6.855 $Y2=1.18
r209 60 62 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.35 $Y=0.415
+ $X2=4.35 $Y2=0.65
r210 56 57 11.0397 $w=5.23e-07 $l=2.25e-07 $layer=LI1_cond $X=2.772 $Y=0.575
+ $X2=2.772 $Y2=0.8
r211 53 56 3.64519 $w=5.23e-07 $l=1.6e-07 $layer=LI1_cond $X=2.772 $Y=0.415
+ $X2=2.772 $Y2=0.575
r212 52 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=1.015
+ $X2=7.335 $Y2=1.18
r213 51 52 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.335 $Y=0.425
+ $X2=7.335 $Y2=1.015
r214 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=2.14 $X2=7.13 $Y2=2.14
r215 46 68 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.13 $Y=1.345
+ $X2=7.13 $Y2=1.18
r216 46 48 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.13 $Y=1.345
+ $X2=7.13 $Y2=2.14
r217 44 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.25 $Y=0.34
+ $X2=7.335 $Y2=0.425
r218 44 45 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=7.25 $Y=0.34
+ $X2=5.65 $Y2=0.34
r219 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.565 $Y=0.425
+ $X2=5.65 $Y2=0.34
r220 42 43 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.565 $Y=0.425
+ $X2=5.565 $Y2=0.565
r221 41 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.65
+ $X2=4.35 $Y2=0.65
r222 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.48 $Y=0.65
+ $X2=5.565 $Y2=0.565
r223 40 41 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=5.48 $Y=0.65
+ $X2=4.435 $Y2=0.65
r224 38 74 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.725
+ $X2=3.33 $Y2=1.89
r225 38 71 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.33 $Y=1.725
+ $X2=3.33 $Y2=1.635
r226 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.33
+ $Y=1.725 $X2=3.33 $Y2=1.725
r227 35 59 4.45426 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=1.725
+ $X2=2.95 $Y2=1.725
r228 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.035 $Y=1.725
+ $X2=3.33 $Y2=1.725
r229 34 53 7.46409 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=3.035 $Y=0.415
+ $X2=2.772 $Y2=0.415
r230 33 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.265 $Y=0.415
+ $X2=4.35 $Y2=0.415
r231 33 34 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.265 $Y=0.415
+ $X2=3.035 $Y2=0.415
r232 32 59 2.3025 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=1.56
+ $X2=2.95 $Y2=1.725
r233 32 57 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.95 $Y=1.56
+ $X2=2.95 $Y2=0.8
r234 27 59 17.036 $w=2.22e-07 $l=3.1e-07 $layer=LI1_cond $X=2.64 $Y=1.725
+ $X2=2.95 $Y2=1.725
r235 27 29 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=2.64 $Y=1.89 $X2=2.64
+ $Y2=1.99
r236 23 49 50.5804 $w=3.46e-07 $l=2.97909e-07 $layer=POLY_cond $X=7.265 $Y=2.39
+ $X2=7.16 $Y2=2.14
r237 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.265 $Y=2.39
+ $X2=7.265 $Y2=2.675
r238 21 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.27
+ $X2=6.855 $Y2=1.27
r239 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.69 $Y=1.27
+ $X2=6.33 $Y2=1.27
r240 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.255 $Y=1.195
+ $X2=6.33 $Y2=1.27
r241 18 20 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.255 $Y=1.195
+ $X2=6.255 $Y2=0.74
r242 14 26 55.5827 $w=2.18e-07 $l=2.62678e-07 $layer=POLY_cond $X=4.005 $Y=1.405
+ $X2=3.935 $Y2=1.635
r243 14 16 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.005 $Y=1.405
+ $X2=4.005 $Y2=0.9
r244 13 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.635
+ $X2=3.33 $Y2=1.635
r245 12 26 11.5617 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.79 $Y=1.635
+ $X2=3.935 $Y2=1.635
r246 12 13 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=3.79 $Y=1.635
+ $X2=3.495 $Y2=1.635
r247 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.4 $Y=2.21 $X2=3.4
+ $Y2=2.495
r248 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.4 $Y=2.12 $X2=3.4
+ $Y2=2.21
r249 8 74 89.4032 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=3.4 $Y=2.12 $X2=3.4
+ $Y2=1.89
r250 2 29 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.83 $X2=2.6 $Y2=1.99
r251 1 56 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.37 $X2=2.675 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%A_830_359# 1 2 7 9 12 16 19 20 25 28 32
c86 16 0 9.2224e-20 $X=4.355 $Y=1.96
c87 12 0 8.87834e-20 $X=4.395 $Y=0.9
r88 31 32 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=6.065 $Y=1.13
+ $X2=6.065 $Y2=1.865
r89 30 31 7.58911 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.985 $Y=0.99
+ $X2=5.985 $Y2=1.13
r90 28 30 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.985 $Y=0.855
+ $X2=5.985 $Y2=0.99
r91 25 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=2.03
+ $X2=6.145 $Y2=1.865
r92 19 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=0.99
+ $X2=5.985 $Y2=0.99
r93 19 20 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=5.82 $Y=0.99
+ $X2=4.445 $Y2=0.99
r94 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.355
+ $Y=1.96 $X2=4.355 $Y2=1.96
r95 14 20 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.355 $Y=1.075
+ $X2=4.445 $Y2=0.99
r96 14 16 54.5303 $w=1.78e-07 $l=8.85e-07 $layer=LI1_cond $X=4.355 $Y=1.075
+ $X2=4.355 $Y2=1.96
r97 10 17 38.6069 $w=3.31e-07 $l=1.92678e-07 $layer=POLY_cond $X=4.395 $Y=1.795
+ $X2=4.335 $Y2=1.96
r98 10 12 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.395 $Y=1.795
+ $X2=4.395 $Y2=0.9
r99 7 17 50.9845 $w=3.31e-07 $l=2.93684e-07 $layer=POLY_cond $X=4.24 $Y=2.21
+ $X2=4.335 $Y2=1.96
r100 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.24 $Y=2.21 $X2=4.24
+ $Y2=2.495
r101 2 25 300 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=1.735 $X2=6.145 $Y2=2.03
r102 1 28 182 $w=1.7e-07 $l=6.8057e-07 $layer=licon1_NDIFF $count=1 $X=5.515
+ $Y=0.37 $X2=5.985 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%A_695_457# 1 2 3 12 14 16 18 19 20 22 23 25
+ 26 30 38 40
c127 38 0 8.87834e-20 $X=4.01 $Y=0.86
r128 36 38 6.67204 $w=3.78e-07 $l=2.2e-07 $layer=LI1_cond $X=3.79 $Y=0.86
+ $X2=4.01 $Y2=0.86
r129 33 34 18.788 $w=2.5e-07 $l=3.85e-07 $layer=LI1_cond $X=3.625 $Y=2.562
+ $X2=4.01 $Y2=2.562
r130 28 40 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.445
+ $X2=4.7 $Y2=2.445
r131 28 30 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=4.785 $Y=2.445
+ $X2=5.085 $Y2=2.445
r132 26 43 72.1174 $w=2.64e-07 $l=3.95e-07 $layer=POLY_cond $X=5.485 $Y=1.452
+ $X2=5.88 $Y2=1.452
r133 26 41 8.21591 $w=2.64e-07 $l=4.5e-08 $layer=POLY_cond $X=5.485 $Y=1.452
+ $X2=5.44 $Y2=1.452
r134 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.485
+ $Y=1.41 $X2=5.485 $Y2=1.41
r135 23 25 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.785 $Y=1.41
+ $X2=5.485 $Y2=1.41
r136 22 40 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.7 $Y=2.32 $X2=4.7
+ $Y2=2.445
r137 21 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.785 $Y2=1.41
r138 21 22 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.7 $Y2=2.32
r139 20 34 5.40474 $w=2.5e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.095 $Y=2.485
+ $X2=4.01 $Y2=2.562
r140 19 40 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.615 $Y=2.485
+ $X2=4.7 $Y2=2.445
r141 19 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.615 $Y=2.485
+ $X2=4.095 $Y2=2.485
r142 18 34 2.99516 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=4.01 $Y=2.4
+ $X2=4.01 $Y2=2.562
r143 17 38 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.01 $Y=1.05
+ $X2=4.01 $Y2=0.86
r144 17 18 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.01 $Y=1.05
+ $X2=4.01 $Y2=2.4
r145 14 43 15.9823 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.88 $Y=1.66
+ $X2=5.88 $Y2=1.452
r146 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.88 $Y=1.66
+ $X2=5.88 $Y2=2.235
r147 10 41 15.9823 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.44 $Y=1.245
+ $X2=5.44 $Y2=1.452
r148 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.44 $Y=1.245
+ $X2=5.44 $Y2=0.74
r149 3 30 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=2.285 $X2=5.085 $Y2=2.485
r150 2 33 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=2.285 $X2=3.625 $Y2=2.52
r151 1 36 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=3.58
+ $Y=0.69 $X2=3.79 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%A_306_74# 1 2 7 9 10 12 14 15 16 17 18 19 21
+ 22 23 24 26 27 32 33 34 37 39 40 44 47 48 52 55 59
c190 55 0 1.09291e-19 $X=1.647 $Y=1.055
c191 52 0 1.65101e-19 $X=2.57 $Y=1.385
c192 14 0 5.68386e-20 $X=2.88 $Y=3.075
r193 61 62 1.78519 $w=4.05e-07 $l=1.5e-08 $layer=POLY_cond $X=2.375 $Y=1.477
+ $X2=2.39 $Y2=1.477
r194 56 59 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.54 $Y=1.975
+ $X2=1.7 $Y2=1.975
r195 53 62 21.4222 $w=4.05e-07 $l=1.8e-07 $layer=POLY_cond $X=2.57 $Y=1.477
+ $X2=2.39 $Y2=1.477
r196 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.385 $X2=2.57 $Y2=1.385
r197 50 52 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=2.57 $Y=1.14
+ $X2=2.57 $Y2=1.385
r198 49 55 3.15366 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.84 $Y=1.055
+ $X2=1.647 $Y2=1.055
r199 48 50 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.57 $Y2=1.14
r200 48 49 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.84 $Y2=1.055
r201 47 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.81
+ $X2=1.54 $Y2=1.975
r202 46 55 3.37808 $w=2.77e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.647 $Y2=1.055
r203 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.54 $Y2=1.81
r204 42 55 3.37808 $w=2.77e-07 $l=8.5e-08 $layer=LI1_cond $X=1.647 $Y=0.97
+ $X2=1.647 $Y2=1.055
r205 42 44 13.6198 $w=3.83e-07 $l=4.55e-07 $layer=LI1_cond $X=1.647 $Y=0.97
+ $X2=1.647 $Y2=0.515
r206 35 37 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.305 $Y=1.585
+ $X2=7.305 $Y2=0.615
r207 33 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.23 $Y=1.66
+ $X2=7.305 $Y2=1.585
r208 33 34 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=7.23 $Y=1.66
+ $X2=6.475 $Y2=1.66
r209 30 40 76.0046 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=6.385 $Y=2.96
+ $X2=6.385 $Y2=3.15
r210 30 32 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.385 $Y=2.96
+ $X2=6.385 $Y2=2.385
r211 29 34 26.9307 $w=1.5e-07 $l=1.89737e-07 $layer=POLY_cond $X=6.385 $Y=1.81
+ $X2=6.475 $Y2=1.66
r212 29 32 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.385 $Y=1.81
+ $X2=6.385 $Y2=2.385
r213 28 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.94 $Y=3.15 $X2=3.85
+ $Y2=3.15
r214 27 40 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.295 $Y=3.15
+ $X2=6.385 $Y2=3.15
r215 27 28 1207.56 $w=1.5e-07 $l=2.355e-06 $layer=POLY_cond $X=6.295 $Y=3.15
+ $X2=3.94 $Y2=3.15
r216 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.85 $Y=2.78
+ $X2=3.85 $Y2=2.495
r217 23 39 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.85 $Y=3.075
+ $X2=3.85 $Y2=3.15
r218 22 24 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.85 $Y=2.87 $X2=3.85
+ $Y2=2.78
r219 22 23 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.85 $Y=2.87
+ $X2=3.85 $Y2=3.075
r220 19 21 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.505 $Y=1.2 $X2=3.505
+ $Y2=0.9
r221 17 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.76 $Y=3.15 $X2=3.85
+ $Y2=3.15
r222 17 18 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.76 $Y=3.15
+ $X2=2.955 $Y2=3.15
r223 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.43 $Y=1.275
+ $X2=3.505 $Y2=1.2
r224 15 16 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=3.43 $Y=1.275
+ $X2=2.955 $Y2=1.275
r225 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.88 $Y=3.075
+ $X2=2.955 $Y2=3.15
r226 13 16 28.9736 $w=4.05e-07 $l=2.36546e-07 $layer=POLY_cond $X=2.88 $Y=1.477
+ $X2=2.955 $Y2=1.275
r227 13 53 36.8938 $w=4.05e-07 $l=3.1e-07 $layer=POLY_cond $X=2.88 $Y=1.477
+ $X2=2.57 $Y2=1.477
r228 13 14 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=2.88 $Y=1.55
+ $X2=2.88 $Y2=3.075
r229 10 62 26.1659 $w=1.5e-07 $l=2.77e-07 $layer=POLY_cond $X=2.39 $Y=1.2
+ $X2=2.39 $Y2=1.477
r230 10 12 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.39 $Y=1.2
+ $X2=2.39 $Y2=0.74
r231 7 61 26.1659 $w=1.5e-07 $l=2.78e-07 $layer=POLY_cond $X=2.375 $Y=1.755
+ $X2=2.375 $Y2=1.477
r232 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.755
+ $X2=2.375 $Y2=2.39
r233 2 59 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.83 $X2=1.7 $Y2=1.975
r234 1 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.53
+ $Y=0.37 $X2=1.675 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%A_1518_203# 1 2 9 10 11 13 16 18 19 25 27 28
+ 30 31 35 38 39 42
r119 38 39 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=8.502 $Y=2.675
+ $X2=8.502 $Y2=2.445
r120 35 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.18
+ $X2=7.755 $Y2=1.345
r121 35 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.18
+ $X2=7.755 $Y2=1.015
r122 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.755
+ $Y=1.18 $X2=7.755 $Y2=1.18
r123 31 34 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.755 $Y=1.1 $X2=7.755
+ $Y2=1.18
r124 29 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.105 $Y=1.185
+ $X2=9.105 $Y2=1.1
r125 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.105 $Y=1.185
+ $X2=9.105 $Y2=1.855
r126 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.02 $Y=1.94
+ $X2=9.105 $Y2=1.855
r127 27 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.02 $Y=1.94
+ $X2=8.685 $Y2=1.94
r128 23 42 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.78 $Y=1.1
+ $X2=9.105 $Y2=1.1
r129 23 25 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=8.78 $Y=1.015 $X2=8.78
+ $Y2=0.615
r130 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.6 $Y=2.025
+ $X2=8.685 $Y2=1.94
r131 21 39 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=8.6 $Y=2.025
+ $X2=8.6 $Y2=2.445
r132 20 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.92 $Y=1.1
+ $X2=7.755 $Y2=1.1
r133 19 23 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=1.1
+ $X2=8.78 $Y2=1.1
r134 19 20 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.615 $Y=1.1
+ $X2=7.92 $Y2=1.1
r135 18 46 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.67 $Y=1.745
+ $X2=7.67 $Y2=1.345
r136 16 45 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.695 $Y=0.615
+ $X2=7.695 $Y2=1.015
r137 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.685 $Y=2.39
+ $X2=7.685 $Y2=2.675
r138 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.685 $Y=2.3
+ $X2=7.685 $Y2=2.39
r139 9 18 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.685 $Y=1.835
+ $X2=7.685 $Y2=1.745
r140 9 10 180.75 $w=1.8e-07 $l=4.65e-07 $layer=POLY_cond $X=7.685 $Y=1.835
+ $X2=7.685 $Y2=2.3
r141 2 38 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=2.465 $X2=8.485 $Y2=2.675
r142 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.64
+ $Y=0.405 $X2=8.78 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%A_1266_74# 1 2 9 12 13 15 16 17 19 21 22 24
+ 25 26 27 29 30 31 32 34 37 39 40 44 45 46 51 54
c161 51 0 1.44605e-19 $X=6.565 $Y=1.6
c162 46 0 1.4888e-19 $X=7.635 $Y=1.6
c163 45 0 3.23044e-20 $X=8.52 $Y=1.6
c164 44 0 1.01622e-19 $X=7.55 $Y=2.475
r165 55 61 3.86218 $w=3.12e-07 $l=2.5e-08 $layer=POLY_cond $X=8.685 $Y=1.52
+ $X2=8.71 $Y2=1.52
r166 55 59 18.5385 $w=3.12e-07 $l=1.2e-07 $layer=POLY_cond $X=8.685 $Y=1.52
+ $X2=8.565 $Y2=1.52
r167 54 57 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.685 $Y=1.52
+ $X2=8.685 $Y2=1.6
r168 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.685
+ $Y=1.52 $X2=8.685 $Y2=1.52
r169 49 51 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.405 $Y=1.6
+ $X2=6.565 $Y2=1.6
r170 45 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.52 $Y=1.6
+ $X2=8.685 $Y2=1.6
r171 45 46 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=8.52 $Y=1.6
+ $X2=7.635 $Y2=1.6
r172 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.55 $Y=1.685
+ $X2=7.635 $Y2=1.6
r173 43 44 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=7.55 $Y=1.685
+ $X2=7.55 $Y2=2.475
r174 40 42 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.65 $Y=2.64
+ $X2=7.04 $Y2=2.64
r175 39 44 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.465 $Y=2.64
+ $X2=7.55 $Y2=2.475
r176 39 42 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.465 $Y=2.64
+ $X2=7.04 $Y2=2.64
r177 35 48 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=0.72
+ $X2=6.405 $Y2=0.72
r178 35 37 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=6.49 $Y=0.72
+ $X2=6.915 $Y2=0.72
r179 34 40 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.565 $Y=2.475
+ $X2=6.65 $Y2=2.64
r180 33 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.565 $Y=1.685
+ $X2=6.565 $Y2=1.6
r181 33 34 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.565 $Y=1.685
+ $X2=6.565 $Y2=2.475
r182 32 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=1.515
+ $X2=6.405 $Y2=1.6
r183 31 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=0.845
+ $X2=6.405 $Y2=0.72
r184 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.405 $Y=0.845
+ $X2=6.405 $Y2=1.515
r185 27 29 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.555 $Y=0.995
+ $X2=9.555 $Y2=0.645
r186 25 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.48 $Y=1.07
+ $X2=9.555 $Y2=0.995
r187 25 26 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=9.48 $Y=1.07
+ $X2=9.305 $Y2=1.07
r188 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.245 $Y=1.97
+ $X2=9.245 $Y2=2.465
r189 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.245 $Y=1.88
+ $X2=9.245 $Y2=1.97
r190 20 30 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.245 $Y=1.685
+ $X2=9.245 $Y2=1.52
r191 20 21 75.7984 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=9.245 $Y=1.685
+ $X2=9.245 $Y2=1.88
r192 19 30 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=9.23 $Y=1.355
+ $X2=9.245 $Y2=1.52
r193 18 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.23 $Y=1.145
+ $X2=9.305 $Y2=1.07
r194 18 19 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.23 $Y=1.145
+ $X2=9.23 $Y2=1.355
r195 17 61 13.3422 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.8 $Y=1.52 $X2=8.71
+ $Y2=1.52
r196 16 30 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.155 $Y=1.52
+ $X2=9.245 $Y2=1.52
r197 16 17 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=9.155 $Y=1.52
+ $X2=8.8 $Y2=1.52
r198 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.71 $Y=2.39
+ $X2=8.71 $Y2=2.675
r199 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.71 $Y=2.3 $X2=8.71
+ $Y2=2.39
r200 11 61 15.628 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.71 $Y=1.685
+ $X2=8.71 $Y2=1.52
r201 11 12 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=8.71 $Y=1.685
+ $X2=8.71 $Y2=2.3
r202 7 59 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.355
+ $X2=8.565 $Y2=1.52
r203 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.565 $Y=1.355
+ $X2=8.565 $Y2=0.615
r204 2 42 300 $w=1.7e-07 $l=1.00395e-06 $layer=licon1_PDIFF $count=2 $X=6.46
+ $Y=1.885 $X2=7.04 $Y2=2.64
r205 1 48 182 $w=1.7e-07 $l=3.79671e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.37 $X2=6.485 $Y2=0.68
r206 1 37 182 $w=1.7e-07 $l=7.23585e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.37 $X2=6.915 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%A_1864_409# 1 2 7 9 12 14 15 18 22 27
r54 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.77
+ $Y=1.55 $X2=9.77 $Y2=1.55
r55 24 27 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=9.47 $Y=1.55 $X2=9.77
+ $Y2=1.55
r56 20 27 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.77 $Y=1.385
+ $X2=9.77 $Y2=1.55
r57 20 22 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=9.77 $Y=1.385
+ $X2=9.77 $Y2=0.645
r58 16 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.47 $Y=1.715
+ $X2=9.47 $Y2=1.55
r59 16 18 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=9.47 $Y=1.715
+ $X2=9.47 $Y2=2.19
r60 14 28 117.157 $w=3.3e-07 $l=6.7e-07 $layer=POLY_cond $X=10.44 $Y=1.55
+ $X2=9.77 $Y2=1.55
r61 14 15 5.03009 $w=3.3e-07 $l=1.01735e-07 $layer=POLY_cond $X=10.44 $Y=1.55
+ $X2=10.53 $Y2=1.575
r62 10 15 37.0704 $w=1.5e-07 $l=1.97358e-07 $layer=POLY_cond $X=10.545 $Y=1.385
+ $X2=10.53 $Y2=1.575
r63 10 12 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=10.545 $Y=1.385
+ $X2=10.545 $Y2=0.74
r64 7 15 37.0704 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=1.575
r65 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=2.4
r66 2 18 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.32
+ $Y=2.045 $X2=9.47 $Y2=2.19
r67 1 22 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.63
+ $Y=0.37 $X2=9.77 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 41 45 51
+ 53 57 59 61 65 67 72 77 85 93 105 108 111 114 117 120 124
r140 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r141 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r142 118 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r143 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r144 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r145 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r146 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r147 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r148 100 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r149 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r150 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r151 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r152 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r153 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r154 94 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=9.02 $Y2=3.33
r155 94 96 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=9.36 $Y2=3.33
r156 93 123 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.595 $Y=3.33
+ $X2=10.817 $Y2=3.33
r157 93 99 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=3.33
+ $X2=10.32 $Y2=3.33
r158 92 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r159 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r160 89 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r161 88 91 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r162 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r163 86 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=3.33
+ $X2=5.645 $Y2=3.33
r164 86 88 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.81 $Y=3.33 $X2=6
+ $Y2=3.33
r165 85 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.805 $Y=3.33
+ $X2=7.97 $Y2=3.33
r166 85 91 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.805 $Y=3.33
+ $X2=7.44 $Y2=3.33
r167 84 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r168 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r169 81 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r170 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r171 80 83 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r172 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r173 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.15 $Y2=3.33
r174 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r175 77 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=3.33
+ $X2=4.55 $Y2=3.33
r176 77 83 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.385 $Y=3.33
+ $X2=4.08 $Y2=3.33
r177 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r178 76 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r179 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r180 73 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.21 $Y2=3.33
r181 73 75 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r182 72 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.15 $Y2=3.33
r183 72 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r184 71 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r185 71 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r186 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r187 68 102 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r188 68 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r189 67 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.21 $Y2=3.33
r190 67 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.72 $Y2=3.33
r191 65 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r192 65 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r193 65 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r194 61 64 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.76 $Y=1.985
+ $X2=10.76 $Y2=2.815
r195 59 123 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.817 $Y2=3.33
r196 59 64 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.76 $Y2=2.815
r197 55 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.02 $Y=3.245
+ $X2=9.02 $Y2=3.33
r198 55 57 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=9.02 $Y=3.245
+ $X2=9.02 $Y2=2.36
r199 54 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.135 $Y=3.33
+ $X2=7.97 $Y2=3.33
r200 53 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.855 $Y=3.33
+ $X2=9.02 $Y2=3.33
r201 53 54 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=8.855 $Y=3.33
+ $X2=8.135 $Y2=3.33
r202 49 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=3.33
r203 49 51 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=2.675
r204 45 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.645 $Y=1.91
+ $X2=5.645 $Y2=2.59
r205 43 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=3.33
r206 43 48 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=2.59
r207 42 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=3.33
+ $X2=4.55 $Y2=3.33
r208 41 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=5.645 $Y2=3.33
r209 41 42 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=4.715 $Y2=3.33
r210 37 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=3.33
r211 37 39 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=2.825
r212 33 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r213 33 35 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.785
r214 29 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.21 $Y2=3.33
r215 29 31 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.21 $Y2=2.815
r216 25 102 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r217 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.23 $Y2=2.75
r218 8 64 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.76 $Y2=2.815
r219 8 61 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.76 $Y2=1.985
r220 7 57 300 $w=1.7e-07 $l=2.82666e-07 $layer=licon1_PDIFF $count=2 $X=8.785
+ $Y=2.465 $X2=9.02 $Y2=2.36
r221 6 51 600 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.465 $X2=7.97 $Y2=2.675
r222 5 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=1.735 $X2=5.645 $Y2=2.59
r223 5 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=1.735 $X2=5.645 $Y2=1.91
r224 4 39 600 $w=1.7e-07 $l=6.46916e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=2.285 $X2=4.55 $Y2=2.825
r225 3 35 600 $w=1.7e-07 $l=1.02727e-06 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.83 $X2=2.15 $Y2=2.785
r226 2 31 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=2.54 $X2=1.17 $Y2=2.815
r227 1 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.27 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%A_30_78# 1 2 3 4 13 16 19 23 25 28 30 34 37
+ 38 39 47
c120 28 0 1.57755e-19 $X=3.67 $Y=2.06
r121 41 43 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=3.135 $Y=2.425
+ $X2=3.135 $Y2=2.495
r122 39 41 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.135 $Y=2.145
+ $X2=3.135 $Y2=2.425
r123 37 38 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.505 $Y=2.41
+ $X2=1.675 $Y2=2.41
r124 34 36 14.9862 $w=2.89e-07 $l=3.55e-07 $layer=LI1_cond $X=0.72 $Y=2.395
+ $X2=0.72 $Y2=2.75
r125 30 32 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.295 $Y=0.6
+ $X2=0.295 $Y2=0.745
r126 27 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=1.39
+ $X2=3.67 $Y2=1.305
r127 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.67 $Y=1.39
+ $X2=3.67 $Y2=2.06
r128 26 39 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.26 $Y=2.145
+ $X2=3.135 $Y2=2.145
r129 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.585 $Y=2.145
+ $X2=3.67 $Y2=2.06
r130 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.585 $Y=2.145
+ $X2=3.26 $Y2=2.145
r131 21 47 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.33 $Y=1.305
+ $X2=3.67 $Y2=1.305
r132 21 23 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=3.33 $Y=1.22
+ $X2=3.33 $Y2=0.9
r133 19 41 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.01 $Y=2.425
+ $X2=3.135 $Y2=2.425
r134 19 38 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=3.01 $Y=2.425
+ $X2=1.675 $Y2=2.425
r135 18 34 3.84173 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=2.395
+ $X2=0.72 $Y2=2.395
r136 18 37 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=0.885 $Y=2.395
+ $X2=1.505 $Y2=2.395
r137 16 34 5.63966 $w=2.89e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.77 $Y=2.31
+ $X2=0.72 $Y2=2.395
r138 15 16 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.77 $Y=0.83
+ $X2=0.77 $Y2=2.31
r139 14 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=0.745
+ $X2=0.295 $Y2=0.745
r140 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.77 $Y2=0.83
r141 13 14 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.46 $Y2=0.745
r142 4 43 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=2.285 $X2=3.175 $Y2=2.495
r143 3 36 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.54 $X2=0.72 $Y2=2.75
r144 2 23 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.69 $X2=3.29 $Y2=0.9
r145 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.39 $X2=0.295 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%Q 1 2 9 13 14 15 16 29
r29 20 32 3.16106 $w=6.98e-07 $l=1.85e-07 $layer=LI1_cond $X=10.075 $Y=2.235
+ $X2=10.075 $Y2=2.05
r30 16 26 0.683473 $w=6.98e-07 $l=4e-08 $layer=LI1_cond $X=10.075 $Y=2.775
+ $X2=10.075 $Y2=2.815
r31 15 16 6.32213 $w=6.98e-07 $l=3.7e-07 $layer=LI1_cond $X=10.075 $Y=2.405
+ $X2=10.075 $Y2=2.775
r32 15 20 2.90476 $w=6.98e-07 $l=1.7e-07 $layer=LI1_cond $X=10.075 $Y=2.405
+ $X2=10.075 $Y2=2.235
r33 14 32 0.256303 $w=6.98e-07 $l=1.5e-08 $layer=LI1_cond $X=10.075 $Y=2.035
+ $X2=10.075 $Y2=2.05
r34 14 29 7.51816 $w=6.98e-07 $l=1.5e-07 $layer=LI1_cond $X=10.075 $Y=2.035
+ $X2=10.075 $Y2=1.885
r35 13 29 33.4652 $w=2.58e-07 $l=7.55e-07 $layer=LI1_cond $X=10.295 $Y=1.13
+ $X2=10.295 $Y2=1.885
r36 7 13 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.33 $Y=0.965
+ $X2=10.33 $Y2=1.13
r37 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=10.33 $Y=0.965
+ $X2=10.33 $Y2=0.515
r38 2 32 400 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.84 $X2=10.26 $Y2=2.05
r39 2 26 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.84 $X2=10.26 $Y2=2.815
r40 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.185
+ $Y=0.37 $X2=10.33 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_1%VGND 1 2 3 4 5 6 21 25 29 33 35 37 40 41 42
+ 48 52 60 68 73 79 89 92 96
c104 29 0 3.23044e-20 $X=7.91 $Y=0.615
r105 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r106 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r107 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r108 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r109 77 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r110 77 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.36 $Y2=0
r111 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r112 74 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.425 $Y=0 $X2=9.3
+ $Y2=0
r113 74 76 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=9.425 $Y=0
+ $X2=10.32 $Y2=0
r114 73 95 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.857 $Y2=0
r115 73 76 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.32 $Y2=0
r116 72 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r117 72 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=7.92
+ $Y2=0
r118 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r119 69 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=7.91
+ $Y2=0
r120 69 71 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=8.075 $Y=0
+ $X2=8.88 $Y2=0
r121 68 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.3
+ $Y2=0
r122 68 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=8.88
+ $Y2=0
r123 67 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r124 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r125 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r126 61 63 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.31 $Y=0 $X2=5.52
+ $Y2=0
r127 60 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.91
+ $Y2=0
r128 60 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r129 59 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r130 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r131 56 59 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r132 56 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r133 55 58 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r134 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r135 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.175
+ $Y2=0
r136 53 55 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.64
+ $Y2=0
r137 52 86 9.04449 $w=3.93e-07 $l=3.1e-07 $layer=LI1_cond $X=5.112 $Y=0
+ $X2=5.112 $Y2=0.31
r138 52 61 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=5.112 $Y=0 $X2=5.31
+ $Y2=0
r139 52 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r140 52 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=4.56 $Y2=0
r141 51 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r142 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r143 48 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.175
+ $Y2=0
r144 48 50 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.68
+ $Y2=0
r145 46 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r146 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r147 42 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=7.44 $Y2=0
r148 42 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r149 42 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r150 40 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r151 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.155
+ $Y2=0
r152 39 50 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r153 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.155
+ $Y2=0
r154 35 95 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.857 $Y2=0
r155 35 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.8 $Y2=0.515
r156 31 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=0.085
+ $X2=9.3 $Y2=0
r157 31 33 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=9.3 $Y=0.085
+ $X2=9.3 $Y2=0.595
r158 27 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r159 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.615
r160 23 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0
r161 23 25 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0.575
r162 19 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r163 19 21 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.6
r164 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.37 $X2=10.76 $Y2=0.515
r165 5 33 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=9.195
+ $Y=0.37 $X2=9.34 $Y2=0.595
r166 4 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.77
+ $Y=0.405 $X2=7.91 $Y2=0.615
r167 3 86 182 $w=1.7e-07 $l=4.89285e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.69 $X2=5.11 $Y2=0.31
r168 2 25 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.37 $X2=2.175 $Y2=0.575
r169 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.39 $X2=1.115 $Y2=0.6
.ends

