* File: sky130_fd_sc_hs__a22oi_2.spice
* Created: Thu Aug 27 20:27:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a22oi_2.pex.spice"
.subckt sky130_fd_sc_hs__a22oi_2  VNB VPB A1 A2 B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_A1_M1003_g N_A_148_74#_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1002 N_A_148_74#_M1003_s N_A2_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_148_74#_M1006_d N_A2_M1006_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1014_d N_A1_M1014_g N_A_148_74#_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.1036 PD=1.28 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1008 N_A_558_74#_M1008_d N_B1_M1008_g N_Y_M1014_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1998 PD=1.13 PS=1.28 NRD=11.34 NRS=25.128 M=1 R=4.93333
+ SA=75002.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_B2_M1013_g N_A_558_74#_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1443 PD=1.02 PS=1.13 NRD=0 NRS=6.48 M=1 R=4.93333 SA=75002.8
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1013_d N_B2_M1015_g N_A_558_74#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1012 N_A_558_74#_M1015_s N_B1_M1012_g N_Y_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_66_368#_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.7 A=0.168 P=2.54 MULT=1
MM1007 N_A_66_368#_M1007_d N_A2_M1007_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_66_368#_M1007_d N_A2_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3416 PD=1.42 PS=1.73 NRD=1.7533 NRS=29.0181 M=1 R=7.46667
+ SA=75001.1 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1009_s N_A1_M1010_g N_A_66_368#_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3416 AS=0.168 PD=1.73 PS=1.42 NRD=29.0181 NRS=1.7533 M=1 R=7.46667
+ SA=75001.9 SB=75002 A=0.168 P=2.54 MULT=1
MM1004 N_A_66_368#_M1010_s N_B1_M1004_g N_Y_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1848 PD=1.42 PS=1.45 NRD=1.7533 NRS=4.3931 M=1 R=7.46667
+ SA=75002.3 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1000 N_A_66_368#_M1000_d N_B2_M1000_g N_Y_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1848 PD=1.42 PS=1.45 NRD=1.7533 NRS=4.3931 M=1 R=7.46667
+ SA=75002.8 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1001 N_A_66_368#_M1000_d N_B2_M1001_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1011 N_A_66_368#_M1011_d N_B1_M1011_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_hs__a22oi_2.pxi.spice"
*
.ends
*
*
