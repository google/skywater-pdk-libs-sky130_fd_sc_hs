* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_126_112# A1_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=8.322e+11p ps=6.72e+06u
M1001 a_117_392# A1_N VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.4e+11p pd=2.48e+06u as=6.446e+11p ps=5.45e+06u
M1002 Y a_126_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 VGND B1 a_488_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1004 a_126_112# A2_N a_117_392# VPB pshort w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1005 a_488_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_399_368# a_126_112# Y VPB pshort w=1.12e+06u l=150000u
+  ad=6.44e+11p pd=5.63e+06u as=3.08e+11p ps=2.79e+06u
M1007 a_399_368# B1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B2 a_399_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2_N a_126_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
