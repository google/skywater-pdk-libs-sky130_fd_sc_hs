* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
X0 VPWR a_922_72# a_340_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_115_74# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 Y A1 a_340_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 a_340_368# a_922_72# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 a_340_368# A1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X5 a_118_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X6 VPWR S a_922_72# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 a_337_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND S a_337_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND a_922_72# a_115_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y A1 a_337_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 Y A0 a_118_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X12 VGND S a_922_72# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_337_74# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR S a_118_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X15 Y A0 a_115_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_115_74# a_922_72# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_118_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
.ends
