* File: sky130_fd_sc_hs__a41o_4.pxi.spice
* Created: Tue Sep  1 19:54:11 2020
* 
x_PM_SKY130_FD_SC_HS__A41O_4%B1 N_B1_M1012_g N_B1_c_139_n N_B1_M1006_g
+ N_B1_M1017_g N_B1_c_140_n N_B1_M1010_g B1 N_B1_c_137_n N_B1_c_138_n
+ PM_SKY130_FD_SC_HS__A41O_4%B1
x_PM_SKY130_FD_SC_HS__A41O_4%A_113_98# N_A_113_98#_M1012_d N_A_113_98#_M1013_d
+ N_A_113_98#_M1006_s N_A_113_98#_c_181_n N_A_113_98#_M1002_g
+ N_A_113_98#_c_182_n N_A_113_98#_M1009_g N_A_113_98#_c_193_n
+ N_A_113_98#_M1000_g N_A_113_98#_c_194_n N_A_113_98#_M1001_g
+ N_A_113_98#_c_183_n N_A_113_98#_M1016_g N_A_113_98#_c_195_n
+ N_A_113_98#_M1003_g N_A_113_98#_c_184_n N_A_113_98#_M1023_g
+ N_A_113_98#_c_196_n N_A_113_98#_M1027_g N_A_113_98#_c_197_n
+ N_A_113_98#_c_230_p N_A_113_98#_c_185_n N_A_113_98#_c_186_n
+ N_A_113_98#_c_187_n N_A_113_98#_c_188_n N_A_113_98#_c_189_n
+ N_A_113_98#_c_190_n N_A_113_98#_c_200_n N_A_113_98#_c_191_n
+ N_A_113_98#_c_192_n PM_SKY130_FD_SC_HS__A41O_4%A_113_98#
x_PM_SKY130_FD_SC_HS__A41O_4%A1 N_A1_c_331_n N_A1_M1005_g N_A1_M1013_g
+ N_A1_c_332_n N_A1_M1008_g N_A1_M1014_g A1 A1 N_A1_c_330_n
+ PM_SKY130_FD_SC_HS__A41O_4%A1
x_PM_SKY130_FD_SC_HS__A41O_4%A2 N_A2_M1011_g N_A2_c_388_n N_A2_M1024_g
+ N_A2_M1026_g N_A2_c_389_n N_A2_M1025_g A2 A2 N_A2_c_387_n
+ PM_SKY130_FD_SC_HS__A41O_4%A2
x_PM_SKY130_FD_SC_HS__A41O_4%A3 N_A3_c_442_n N_A3_M1019_g N_A3_M1007_g
+ N_A3_c_443_n N_A3_M1021_g N_A3_M1018_g A3 A3 A3 N_A3_c_441_n
+ PM_SKY130_FD_SC_HS__A41O_4%A3
x_PM_SKY130_FD_SC_HS__A41O_4%A4 N_A4_c_500_n N_A4_M1020_g N_A4_M1004_g
+ N_A4_c_501_n N_A4_M1022_g N_A4_M1015_g A4 A4 N_A4_c_499_n
+ PM_SKY130_FD_SC_HS__A41O_4%A4
x_PM_SKY130_FD_SC_HS__A41O_4%A_27_392# N_A_27_392#_M1006_d N_A_27_392#_M1010_d
+ N_A_27_392#_M1005_s N_A_27_392#_M1024_d N_A_27_392#_M1019_s
+ N_A_27_392#_M1020_d N_A_27_392#_c_537_n N_A_27_392#_c_538_n
+ N_A_27_392#_c_539_n N_A_27_392#_c_540_n N_A_27_392#_c_541_n
+ N_A_27_392#_c_542_n N_A_27_392#_c_543_n N_A_27_392#_c_588_n
+ N_A_27_392#_c_544_n N_A_27_392#_c_545_n N_A_27_392#_c_546_n
+ N_A_27_392#_c_547_n N_A_27_392#_c_548_n N_A_27_392#_c_549_n
+ N_A_27_392#_c_550_n N_A_27_392#_c_565_n N_A_27_392#_c_551_n
+ N_A_27_392#_c_552_n N_A_27_392#_c_553_n PM_SKY130_FD_SC_HS__A41O_4%A_27_392#
x_PM_SKY130_FD_SC_HS__A41O_4%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1027_d
+ N_VPWR_M1008_d N_VPWR_M1025_s N_VPWR_M1021_d N_VPWR_M1022_s N_VPWR_c_673_n
+ N_VPWR_c_674_n N_VPWR_c_675_n N_VPWR_c_676_n N_VPWR_c_677_n N_VPWR_c_678_n
+ N_VPWR_c_679_n N_VPWR_c_680_n N_VPWR_c_681_n N_VPWR_c_682_n VPWR
+ N_VPWR_c_683_n N_VPWR_c_684_n N_VPWR_c_685_n N_VPWR_c_686_n N_VPWR_c_687_n
+ N_VPWR_c_688_n N_VPWR_c_689_n N_VPWR_c_690_n N_VPWR_c_691_n N_VPWR_c_692_n
+ N_VPWR_c_693_n N_VPWR_c_672_n PM_SKY130_FD_SC_HS__A41O_4%VPWR
x_PM_SKY130_FD_SC_HS__A41O_4%X N_X_M1002_s N_X_M1016_s N_X_M1000_s N_X_M1003_s
+ N_X_c_783_n N_X_c_790_n N_X_c_794_n X X X N_X_c_805_n
+ PM_SKY130_FD_SC_HS__A41O_4%X
x_PM_SKY130_FD_SC_HS__A41O_4%VGND N_VGND_M1012_s N_VGND_M1017_s N_VGND_M1009_d
+ N_VGND_M1023_d N_VGND_M1004_s N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n
+ N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n VGND
+ N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n
+ N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n
+ PM_SKY130_FD_SC_HS__A41O_4%VGND
x_PM_SKY130_FD_SC_HS__A41O_4%A_751_74# N_A_751_74#_M1013_s N_A_751_74#_M1014_s
+ N_A_751_74#_M1026_d N_A_751_74#_c_917_n N_A_751_74#_c_918_n
+ N_A_751_74#_c_919_n N_A_751_74#_c_920_n N_A_751_74#_c_921_n
+ N_A_751_74#_c_922_n PM_SKY130_FD_SC_HS__A41O_4%A_751_74#
x_PM_SKY130_FD_SC_HS__A41O_4%A_1010_74# N_A_1010_74#_M1011_s
+ N_A_1010_74#_M1007_s N_A_1010_74#_c_960_n N_A_1010_74#_c_957_n
+ N_A_1010_74#_c_958_n N_A_1010_74#_c_979_p
+ PM_SKY130_FD_SC_HS__A41O_4%A_1010_74#
x_PM_SKY130_FD_SC_HS__A41O_4%A_1205_74# N_A_1205_74#_M1007_d
+ N_A_1205_74#_M1018_d N_A_1205_74#_M1015_d N_A_1205_74#_c_981_n
+ N_A_1205_74#_c_982_n N_A_1205_74#_c_983_n N_A_1205_74#_c_993_n
+ N_A_1205_74#_c_984_n N_A_1205_74#_c_985_n N_A_1205_74#_c_986_n
+ PM_SKY130_FD_SC_HS__A41O_4%A_1205_74#
cc_1 VNB N_B1_M1012_g 0.028167f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.86
cc_2 VNB N_B1_M1017_g 0.0217362f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.86
cc_3 VNB N_B1_c_137_n 0.00897124f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_4 VNB N_B1_c_138_n 0.0399762f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.667
cc_5 VNB N_A_113_98#_c_181_n 0.0178666f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.86
cc_6 VNB N_A_113_98#_c_182_n 0.0175516f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.46
cc_7 VNB N_A_113_98#_c_183_n 0.0170902f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.667
cc_8 VNB N_A_113_98#_c_184_n 0.0175501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_113_98#_c_185_n 0.0103055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_113_98#_c_186_n 0.00952083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_113_98#_c_187_n 0.00190145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_113_98#_c_188_n 0.00624434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_113_98#_c_189_n 0.00766989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_113_98#_c_190_n 0.00374035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_113_98#_c_191_n 0.00201479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_113_98#_c_192_n 0.109327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_M1013_g 0.0371828f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_18 VNB N_A1_M1014_g 0.0287381f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.46
cc_19 VNB A1 0.0104715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_330_n 0.0357649f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_21 VNB N_A2_M1011_g 0.028526f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.86
cc_22 VNB N_A2_M1026_g 0.036548f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.86
cc_23 VNB A2 0.00550923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_387_n 0.0315849f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_25 VNB N_A3_M1007_g 0.0362365f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_26 VNB N_A3_M1018_g 0.0274595f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.46
cc_27 VNB A3 0.00738038f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.667
cc_28 VNB N_A3_c_441_n 0.0314257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A4_M1004_g 0.0272452f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_30 VNB N_A4_M1015_g 0.0376705f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.46
cc_31 VNB A4 0.0120975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A4_c_499_n 0.0274019f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_33 VNB N_VPWR_c_672_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.00448002f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_35 VNB N_VGND_c_820_n 0.0105185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_821_n 0.0526721f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_37 VNB N_VGND_c_822_n 0.0173083f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.667
cc_38 VNB N_VGND_c_823_n 0.0141935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_824_n 0.0184332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_825_n 0.00673507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_826_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_827_n 0.018961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_828_n 0.0187092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_829_n 0.0962806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_830_n 0.0171537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_831_n 0.448983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_832_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_833_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_834_n 0.00477852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_835_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_751_74#_c_917_n 0.0103454f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.86
cc_52 VNB N_A_751_74#_c_918_n 0.00171068f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.885
cc_53 VNB N_A_751_74#_c_919_n 0.00722456f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.46
cc_54 VNB N_A_751_74#_c_920_n 0.00272742f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.46
cc_55 VNB N_A_751_74#_c_921_n 0.0020013f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.667
cc_56 VNB N_A_751_74#_c_922_n 0.00842315f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_57 VNB N_A_1010_74#_c_957_n 0.0296356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1010_74#_c_958_n 0.00186312f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.885
cc_59 VNB N_A_1205_74#_c_981_n 0.00473932f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.885
cc_60 VNB N_A_1205_74#_c_982_n 0.00450918f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.46
cc_61 VNB N_A_1205_74#_c_983_n 0.00471344f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_62 VNB N_A_1205_74#_c_984_n 0.0195741f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.667
cc_63 VNB N_A_1205_74#_c_985_n 0.00239138f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.667
cc_64 VNB N_A_1205_74#_c_986_n 0.0306368f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_65 VPB N_B1_c_139_n 0.0190805f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_66 VPB N_B1_c_140_n 0.0187112f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.885
cc_67 VPB N_B1_c_137_n 0.0054581f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_68 VPB N_B1_c_138_n 0.0557752f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.667
cc_69 VPB N_A_113_98#_c_193_n 0.0190933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_113_98#_c_194_n 0.0150314f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_71 VPB N_A_113_98#_c_195_n 0.0144483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_113_98#_c_196_n 0.0153756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_113_98#_c_197_n 0.00136951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_113_98#_c_185_n 0.00145238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_113_98#_c_187_n 0.00164501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_113_98#_c_200_n 0.00353907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_113_98#_c_192_n 0.0693763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A1_c_331_n 0.0178959f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=1.45
cc_79 VPB N_A1_c_332_n 0.0186451f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.45
cc_80 VPB A1 0.00589024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A1_c_330_n 0.0428573f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_82 VPB N_A2_c_388_n 0.0171687f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_83 VPB N_A2_c_389_n 0.0164749f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.885
cc_84 VPB A2 0.00147646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A2_c_387_n 0.0416008f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_86 VPB N_A3_c_442_n 0.0168629f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=1.45
cc_87 VPB N_A3_c_443_n 0.0158613f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.45
cc_88 VPB A3 0.00576921f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.667
cc_89 VPB N_A3_c_441_n 0.0376793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A4_c_500_n 0.0161547f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=1.45
cc_91 VPB N_A4_c_501_n 0.0179591f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.45
cc_92 VPB A4 0.00947347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A4_c_499_n 0.0371299f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_94 VPB N_A_27_392#_c_537_n 0.0387674f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.667
cc_95 VPB N_A_27_392#_c_538_n 0.0068066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_392#_c_539_n 0.00983167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_392#_c_540_n 0.00876326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_27_392#_c_541_n 0.00500154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_27_392#_c_542_n 0.0127254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_392#_c_543_n 0.00307639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_392#_c_544_n 0.0118851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_392#_c_545_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_392#_c_546_n 0.00469417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_392#_c_547_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_27_392#_c_548_n 0.0033885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_27_392#_c_549_n 0.00201669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_392#_c_550_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_392#_c_551_n 0.00332867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_392#_c_552_n 0.00183558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_392#_c_553_n 0.00193086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_673_n 0.00895772f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_112 VPB N_VPWR_c_674_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_675_n 0.00614032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_676_n 0.0104924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_677_n 0.00830446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_678_n 0.00596713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_679_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_680_n 0.0519123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_681_n 0.024741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_682_n 0.0088221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_683_n 0.041497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_684_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_685_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_686_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_687_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_688_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_689_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_690_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_691_n 0.00652596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_692_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_693_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_672_n 0.115168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB X 0.00180702f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_134 N_B1_M1017_g N_A_113_98#_c_181_n 0.0235643f $X=0.92 $Y=0.86 $X2=0 $Y2=0
cc_135 N_B1_c_139_n N_A_113_98#_c_197_n 0.00420635f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_136 N_B1_c_138_n N_A_113_98#_c_197_n 0.00462586f $X=0.92 $Y=1.667 $X2=0 $Y2=0
cc_137 N_B1_M1012_g N_A_113_98#_c_185_n 0.0164959f $X=0.49 $Y=0.86 $X2=0 $Y2=0
cc_138 N_B1_M1017_g N_A_113_98#_c_185_n 0.0311738f $X=0.92 $Y=0.86 $X2=0 $Y2=0
cc_139 N_B1_c_137_n N_A_113_98#_c_185_n 0.0185991f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_140 N_B1_c_138_n N_A_113_98#_c_185_n 0.0290194f $X=0.92 $Y=1.667 $X2=0 $Y2=0
cc_141 N_B1_c_139_n N_A_113_98#_c_200_n 0.00142223f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_142 N_B1_c_140_n N_A_113_98#_c_200_n 0.00188735f $X=1.005 $Y=1.885 $X2=0
+ $Y2=0
cc_143 N_B1_c_137_n N_A_113_98#_c_200_n 0.00804179f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_144 N_B1_c_138_n N_A_113_98#_c_200_n 0.015845f $X=0.92 $Y=1.667 $X2=0 $Y2=0
cc_145 N_B1_M1017_g N_A_113_98#_c_192_n 0.00330336f $X=0.92 $Y=0.86 $X2=0 $Y2=0
cc_146 N_B1_c_138_n N_A_113_98#_c_192_n 0.0100743f $X=0.92 $Y=1.667 $X2=0 $Y2=0
cc_147 N_B1_c_139_n N_A_27_392#_c_537_n 0.011006f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_148 N_B1_c_140_n N_A_27_392#_c_537_n 6.2649e-19 $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_149 N_B1_c_137_n N_A_27_392#_c_537_n 0.0272312f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_150 N_B1_c_138_n N_A_27_392#_c_537_n 0.00500623f $X=0.92 $Y=1.667 $X2=0 $Y2=0
cc_151 N_B1_c_139_n N_A_27_392#_c_538_n 0.0111147f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_152 N_B1_c_140_n N_A_27_392#_c_538_n 0.013744f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_153 N_B1_c_139_n N_A_27_392#_c_539_n 0.00262934f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_154 N_B1_c_140_n N_A_27_392#_c_540_n 0.00401595f $X=1.005 $Y=1.885 $X2=0
+ $Y2=0
cc_155 N_B1_c_138_n N_A_27_392#_c_540_n 4.54337e-19 $X=0.92 $Y=1.667 $X2=0 $Y2=0
cc_156 N_B1_c_139_n N_A_27_392#_c_541_n 5.79827e-19 $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_157 N_B1_c_140_n N_A_27_392#_c_541_n 0.00578081f $X=1.005 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_B1_c_140_n N_A_27_392#_c_565_n 0.00164802f $X=1.005 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_B1_c_140_n N_VPWR_c_673_n 0.0013297f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_160 N_B1_c_139_n N_VPWR_c_683_n 0.00278257f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_161 N_B1_c_140_n N_VPWR_c_683_n 0.00278257f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_162 N_B1_c_139_n N_VPWR_c_672_n 0.00357777f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_163 N_B1_c_140_n N_VPWR_c_672_n 0.00359084f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_164 N_B1_M1012_g N_VGND_c_821_n 0.00650665f $X=0.49 $Y=0.86 $X2=0 $Y2=0
cc_165 N_B1_c_137_n N_VGND_c_821_n 0.0178692f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_166 N_B1_c_138_n N_VGND_c_821_n 0.00318891f $X=0.92 $Y=1.667 $X2=0 $Y2=0
cc_167 N_B1_M1017_g N_VGND_c_822_n 0.00339639f $X=0.92 $Y=0.86 $X2=0 $Y2=0
cc_168 N_B1_M1012_g N_VGND_c_827_n 0.00472523f $X=0.49 $Y=0.86 $X2=0 $Y2=0
cc_169 N_B1_M1017_g N_VGND_c_827_n 0.00378531f $X=0.92 $Y=0.86 $X2=0 $Y2=0
cc_170 N_B1_M1012_g N_VGND_c_831_n 0.00508379f $X=0.49 $Y=0.86 $X2=0 $Y2=0
cc_171 N_B1_M1017_g N_VGND_c_831_n 0.00508379f $X=0.92 $Y=0.86 $X2=0 $Y2=0
cc_172 N_A_113_98#_c_196_n N_A1_c_331_n 0.0311429f $X=3.365 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_113_98#_c_186_n N_A1_M1013_g 0.00105344f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_174 N_A_113_98#_c_188_n N_A1_M1013_g 0.00461429f $X=3.56 $Y=0.66 $X2=0 $Y2=0
cc_175 N_A_113_98#_c_189_n N_A1_M1013_g 0.00996456f $X=4.165 $Y=0.34 $X2=0 $Y2=0
cc_176 N_A_113_98#_c_191_n N_A1_M1013_g 0.00608359f $X=4.33 $Y=0.34 $X2=0 $Y2=0
cc_177 N_A_113_98#_c_192_n N_A1_M1013_g 0.0032087f $X=2.935 $Y=1.552 $X2=0 $Y2=0
cc_178 N_A_113_98#_c_191_n N_A1_M1014_g 0.00594068f $X=4.33 $Y=0.34 $X2=0 $Y2=0
cc_179 N_A_113_98#_c_186_n A1 0.00565806f $X=3.475 $Y=0.745 $X2=0 $Y2=0
cc_180 N_A_113_98#_c_192_n A1 0.00350993f $X=2.935 $Y=1.552 $X2=0 $Y2=0
cc_181 N_A_113_98#_c_196_n N_A1_c_330_n 0.00424277f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_113_98#_c_192_n N_A1_c_330_n 0.010539f $X=2.935 $Y=1.552 $X2=0 $Y2=0
cc_183 N_A_113_98#_c_191_n N_A2_M1011_g 4.65448e-19 $X=4.33 $Y=0.34 $X2=0 $Y2=0
cc_184 N_A_113_98#_c_197_n N_A_27_392#_c_537_n 0.0298193f $X=0.752 $Y=2.087
+ $X2=0 $Y2=0
cc_185 N_A_113_98#_M1006_s N_A_27_392#_c_538_n 0.00250873f $X=0.58 $Y=1.96 $X2=0
+ $Y2=0
cc_186 N_A_113_98#_c_193_n N_A_27_392#_c_538_n 6.15812e-19 $X=2.015 $Y=1.765
+ $X2=0 $Y2=0
cc_187 N_A_113_98#_c_230_p N_A_27_392#_c_538_n 0.0179627f $X=0.78 $Y=2.115 $X2=0
+ $Y2=0
cc_188 N_A_113_98#_c_193_n N_A_27_392#_c_540_n 0.00876419f $X=2.015 $Y=1.765
+ $X2=0 $Y2=0
cc_189 N_A_113_98#_c_185_n N_A_27_392#_c_540_n 0.0105623f $X=0.805 $Y=1.67 $X2=0
+ $Y2=0
cc_190 N_A_113_98#_c_187_n N_A_27_392#_c_540_n 0.0107097f $X=2.22 $Y=1.505 $X2=0
+ $Y2=0
cc_191 N_A_113_98#_c_200_n N_A_27_392#_c_540_n 0.0134828f $X=0.752 $Y=1.95 $X2=0
+ $Y2=0
cc_192 N_A_113_98#_c_192_n N_A_27_392#_c_540_n 4.18568e-19 $X=2.935 $Y=1.552
+ $X2=0 $Y2=0
cc_193 N_A_113_98#_c_193_n N_A_27_392#_c_541_n 0.00345021f $X=2.015 $Y=1.765
+ $X2=0 $Y2=0
cc_194 N_A_113_98#_c_193_n N_A_27_392#_c_542_n 0.0184914f $X=2.015 $Y=1.765
+ $X2=0 $Y2=0
cc_195 N_A_113_98#_c_194_n N_A_27_392#_c_542_n 0.0146711f $X=2.465 $Y=1.765
+ $X2=0 $Y2=0
cc_196 N_A_113_98#_c_195_n N_A_27_392#_c_542_n 0.0146649f $X=2.915 $Y=1.765
+ $X2=0 $Y2=0
cc_197 N_A_113_98#_c_196_n N_A_27_392#_c_542_n 0.0191001f $X=3.365 $Y=1.765
+ $X2=0 $Y2=0
cc_198 N_A_113_98#_c_187_n N_A_27_392#_c_542_n 0.0173701f $X=2.22 $Y=1.505 $X2=0
+ $Y2=0
cc_199 N_A_113_98#_c_192_n N_A_27_392#_c_542_n 0.0106022f $X=2.935 $Y=1.552
+ $X2=0 $Y2=0
cc_200 N_A_113_98#_c_193_n N_VPWR_c_673_n 0.0113718f $X=2.015 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A_113_98#_c_194_n N_VPWR_c_673_n 0.00136002f $X=2.465 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_113_98#_c_193_n N_VPWR_c_674_n 0.00136002f $X=2.015 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_113_98#_c_194_n N_VPWR_c_674_n 0.0102964f $X=2.465 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A_113_98#_c_195_n N_VPWR_c_674_n 0.0103024f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A_113_98#_c_196_n N_VPWR_c_674_n 0.0013959f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_113_98#_c_195_n N_VPWR_c_675_n 0.0013005f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_113_98#_c_196_n N_VPWR_c_675_n 0.00984264f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_113_98#_c_193_n N_VPWR_c_684_n 0.00413917f $X=2.015 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_113_98#_c_194_n N_VPWR_c_684_n 0.00413917f $X=2.465 $Y=1.765 $X2=0
+ $Y2=0
cc_210 N_A_113_98#_c_195_n N_VPWR_c_685_n 0.00413917f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_A_113_98#_c_196_n N_VPWR_c_685_n 0.00413917f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_A_113_98#_c_193_n N_VPWR_c_672_n 0.00817726f $X=2.015 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A_113_98#_c_194_n N_VPWR_c_672_n 0.00817726f $X=2.465 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A_113_98#_c_195_n N_VPWR_c_672_n 0.00817726f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_A_113_98#_c_196_n N_VPWR_c_672_n 0.00817726f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_216 N_A_113_98#_c_186_n N_X_M1002_s 0.0046269f $X=3.475 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_113_98#_c_186_n N_X_M1016_s 0.00462302f $X=3.475 $Y=0.745 $X2=0 $Y2=0
cc_218 N_A_113_98#_c_181_n N_X_c_783_n 0.00300964f $X=1.5 $Y=1.34 $X2=0 $Y2=0
cc_219 N_A_113_98#_c_182_n N_X_c_783_n 0.0091829f $X=1.93 $Y=1.34 $X2=0 $Y2=0
cc_220 N_A_113_98#_c_183_n N_X_c_783_n 0.0099061f $X=2.505 $Y=1.34 $X2=0 $Y2=0
cc_221 N_A_113_98#_c_185_n N_X_c_783_n 0.00889978f $X=0.805 $Y=1.67 $X2=0 $Y2=0
cc_222 N_A_113_98#_c_186_n N_X_c_783_n 0.0548785f $X=3.475 $Y=0.745 $X2=0 $Y2=0
cc_223 N_A_113_98#_c_187_n N_X_c_783_n 0.0545167f $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_224 N_A_113_98#_c_192_n N_X_c_783_n 0.00774711f $X=2.935 $Y=1.552 $X2=0 $Y2=0
cc_225 N_A_113_98#_c_193_n N_X_c_790_n 0.0132549f $X=2.015 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A_113_98#_c_194_n N_X_c_790_n 0.0137399f $X=2.465 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A_113_98#_c_187_n N_X_c_790_n 0.0194227f $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_228 N_A_113_98#_c_192_n N_X_c_790_n 0.00605684f $X=2.935 $Y=1.552 $X2=0 $Y2=0
cc_229 N_A_113_98#_c_183_n N_X_c_794_n 7.32094e-19 $X=2.505 $Y=1.34 $X2=0 $Y2=0
cc_230 N_A_113_98#_c_184_n N_X_c_794_n 0.00795334f $X=2.935 $Y=1.34 $X2=0 $Y2=0
cc_231 N_A_113_98#_c_186_n N_X_c_794_n 0.0460704f $X=3.475 $Y=0.745 $X2=0 $Y2=0
cc_232 N_A_113_98#_c_182_n X 7.60222e-19 $X=1.93 $Y=1.34 $X2=0 $Y2=0
cc_233 N_A_113_98#_c_194_n X 0.00247845f $X=2.465 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_113_98#_c_183_n X 0.00500527f $X=2.505 $Y=1.34 $X2=0 $Y2=0
cc_235 N_A_113_98#_c_195_n X 0.0027293f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A_113_98#_c_184_n X 0.00702286f $X=2.935 $Y=1.34 $X2=0 $Y2=0
cc_237 N_A_113_98#_c_196_n X 0.00226866f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_113_98#_c_187_n X 0.0276335f $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_239 N_A_113_98#_c_192_n X 0.0649664f $X=2.935 $Y=1.552 $X2=0 $Y2=0
cc_240 N_A_113_98#_c_195_n N_X_c_805_n 0.00963276f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_113_98#_c_196_n N_X_c_805_n 0.00591774f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_113_98#_c_185_n N_VGND_M1017_s 0.00780828f $X=0.805 $Y=1.67 $X2=0
+ $Y2=0
cc_243 N_A_113_98#_c_186_n N_VGND_M1017_s 0.00402935f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_244 N_A_113_98#_c_186_n N_VGND_M1009_d 0.0068273f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_245 N_A_113_98#_c_186_n N_VGND_M1023_d 0.0083134f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_246 N_A_113_98#_c_185_n N_VGND_c_821_n 0.0320582f $X=0.805 $Y=1.67 $X2=0
+ $Y2=0
cc_247 N_A_113_98#_c_181_n N_VGND_c_822_n 0.00379005f $X=1.5 $Y=1.34 $X2=0 $Y2=0
cc_248 N_A_113_98#_c_185_n N_VGND_c_822_n 0.0164999f $X=0.805 $Y=1.67 $X2=0
+ $Y2=0
cc_249 N_A_113_98#_c_186_n N_VGND_c_822_n 0.0112155f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_250 N_A_113_98#_c_182_n N_VGND_c_823_n 0.00378243f $X=1.93 $Y=1.34 $X2=0
+ $Y2=0
cc_251 N_A_113_98#_c_183_n N_VGND_c_823_n 0.0021586f $X=2.505 $Y=1.34 $X2=0
+ $Y2=0
cc_252 N_A_113_98#_c_186_n N_VGND_c_823_n 0.0246365f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_253 N_A_113_98#_c_183_n N_VGND_c_824_n 0.0038134f $X=2.505 $Y=1.34 $X2=0
+ $Y2=0
cc_254 N_A_113_98#_c_184_n N_VGND_c_824_n 0.0038134f $X=2.935 $Y=1.34 $X2=0
+ $Y2=0
cc_255 N_A_113_98#_c_186_n N_VGND_c_824_n 0.00922288f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_256 N_A_113_98#_c_184_n N_VGND_c_825_n 0.00379495f $X=2.935 $Y=1.34 $X2=0
+ $Y2=0
cc_257 N_A_113_98#_c_186_n N_VGND_c_825_n 0.0186889f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_258 N_A_113_98#_c_188_n N_VGND_c_825_n 0.00491052f $X=3.56 $Y=0.66 $X2=0
+ $Y2=0
cc_259 N_A_113_98#_c_190_n N_VGND_c_825_n 0.0145179f $X=3.645 $Y=0.34 $X2=0
+ $Y2=0
cc_260 N_A_113_98#_c_185_n N_VGND_c_827_n 0.0123334f $X=0.805 $Y=1.67 $X2=0
+ $Y2=0
cc_261 N_A_113_98#_c_181_n N_VGND_c_828_n 0.0038134f $X=1.5 $Y=1.34 $X2=0 $Y2=0
cc_262 N_A_113_98#_c_182_n N_VGND_c_828_n 0.0038134f $X=1.93 $Y=1.34 $X2=0 $Y2=0
cc_263 N_A_113_98#_c_186_n N_VGND_c_828_n 0.00931454f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_264 N_A_113_98#_c_186_n N_VGND_c_829_n 0.00287846f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_265 N_A_113_98#_c_189_n N_VGND_c_829_n 0.0331045f $X=4.165 $Y=0.34 $X2=0
+ $Y2=0
cc_266 N_A_113_98#_c_190_n N_VGND_c_829_n 0.0120335f $X=3.645 $Y=0.34 $X2=0
+ $Y2=0
cc_267 N_A_113_98#_c_191_n N_VGND_c_829_n 0.0222074f $X=4.33 $Y=0.34 $X2=0 $Y2=0
cc_268 N_A_113_98#_c_181_n N_VGND_c_831_n 0.00508379f $X=1.5 $Y=1.34 $X2=0 $Y2=0
cc_269 N_A_113_98#_c_182_n N_VGND_c_831_n 0.00508379f $X=1.93 $Y=1.34 $X2=0
+ $Y2=0
cc_270 N_A_113_98#_c_183_n N_VGND_c_831_n 0.00508379f $X=2.505 $Y=1.34 $X2=0
+ $Y2=0
cc_271 N_A_113_98#_c_184_n N_VGND_c_831_n 0.00508379f $X=2.935 $Y=1.34 $X2=0
+ $Y2=0
cc_272 N_A_113_98#_c_185_n N_VGND_c_831_n 0.0171981f $X=0.805 $Y=1.67 $X2=0
+ $Y2=0
cc_273 N_A_113_98#_c_186_n N_VGND_c_831_n 0.0452434f $X=3.475 $Y=0.745 $X2=0
+ $Y2=0
cc_274 N_A_113_98#_c_189_n N_VGND_c_831_n 0.018978f $X=4.165 $Y=0.34 $X2=0 $Y2=0
cc_275 N_A_113_98#_c_190_n N_VGND_c_831_n 0.00658039f $X=3.645 $Y=0.34 $X2=0
+ $Y2=0
cc_276 N_A_113_98#_c_191_n N_VGND_c_831_n 0.0123185f $X=4.33 $Y=0.34 $X2=0 $Y2=0
cc_277 N_A_113_98#_c_189_n N_A_751_74#_M1013_s 0.00482965f $X=4.165 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_278 N_A_113_98#_M1013_d N_A_751_74#_c_917_n 0.00177314f $X=4.19 $Y=0.37 $X2=0
+ $Y2=0
cc_279 N_A_113_98#_c_189_n N_A_751_74#_c_917_n 0.00440398f $X=4.165 $Y=0.34
+ $X2=0 $Y2=0
cc_280 N_A_113_98#_c_191_n N_A_751_74#_c_917_n 0.016611f $X=4.33 $Y=0.34 $X2=0
+ $Y2=0
cc_281 N_A_113_98#_c_191_n N_A_751_74#_c_918_n 0.0114662f $X=4.33 $Y=0.34 $X2=0
+ $Y2=0
cc_282 N_A_113_98#_c_186_n N_A_751_74#_c_921_n 0.0112805f $X=3.475 $Y=0.745
+ $X2=0 $Y2=0
cc_283 N_A_113_98#_c_189_n N_A_751_74#_c_921_n 0.00817883f $X=4.165 $Y=0.34
+ $X2=0 $Y2=0
cc_284 N_A1_M1014_g N_A2_M1011_g 0.020505f $X=4.545 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A1_c_332_n N_A2_c_388_n 0.019526f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_286 N_A1_c_330_n A2 0.00242024f $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_287 N_A1_c_330_n N_A2_c_387_n 0.0237682f $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_288 N_A1_c_331_n N_A_27_392#_c_542_n 0.0176536f $X=3.885 $Y=1.885 $X2=0 $Y2=0
cc_289 A1 N_A_27_392#_c_542_n 0.0164848f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_290 N_A1_c_330_n N_A_27_392#_c_542_n 0.00109095f $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_291 N_A1_c_331_n N_A_27_392#_c_543_n 0.00560351f $X=3.885 $Y=1.885 $X2=0
+ $Y2=0
cc_292 A1 N_A_27_392#_c_543_n 0.01265f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_293 N_A1_c_330_n N_A_27_392#_c_543_n 0.0124207f $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_294 N_A1_c_331_n N_A_27_392#_c_588_n 0.00481222f $X=3.885 $Y=1.885 $X2=0
+ $Y2=0
cc_295 N_A1_c_332_n N_A_27_392#_c_588_n 0.00484336f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_296 N_A1_c_332_n N_A_27_392#_c_544_n 0.0213571f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_297 N_A1_c_330_n N_A_27_392#_c_544_n 0.00405701f $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_298 N_A1_c_332_n N_A_27_392#_c_545_n 8.2453e-19 $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_299 N_A1_c_331_n N_A_27_392#_c_551_n 0.00904308f $X=3.885 $Y=1.885 $X2=0
+ $Y2=0
cc_300 N_A1_c_332_n N_A_27_392#_c_551_n 0.00772304f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_301 N_A1_c_331_n N_VPWR_c_675_n 0.00513483f $X=3.885 $Y=1.885 $X2=0 $Y2=0
cc_302 N_A1_c_332_n N_VPWR_c_676_n 0.0088525f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_303 N_A1_c_331_n N_VPWR_c_681_n 0.00461464f $X=3.885 $Y=1.885 $X2=0 $Y2=0
cc_304 N_A1_c_332_n N_VPWR_c_681_n 0.00461464f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_305 N_A1_c_331_n N_VPWR_c_672_n 0.00910527f $X=3.885 $Y=1.885 $X2=0 $Y2=0
cc_306 N_A1_c_332_n N_VPWR_c_672_n 0.00911487f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_307 A1 X 0.0279316f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_308 N_A1_c_330_n X 4.98655e-19 $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_309 N_A1_c_331_n N_X_c_805_n 0.00107036f $X=3.885 $Y=1.885 $X2=0 $Y2=0
cc_310 N_A1_c_330_n N_X_c_805_n 2.11258e-19 $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_311 N_A1_M1013_g N_VGND_c_829_n 0.00279469f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A1_M1014_g N_VGND_c_829_n 0.0043213f $X=4.545 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A1_M1013_g N_VGND_c_831_n 0.00357517f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A1_M1014_g N_VGND_c_831_n 0.00432202f $X=4.545 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A1_M1013_g N_A_751_74#_c_917_n 0.0171916f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A1_M1014_g N_A_751_74#_c_917_n 0.0208153f $X=4.545 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A1_c_330_n N_A_751_74#_c_917_n 0.00357612f $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_318 N_A1_M1014_g N_A_751_74#_c_918_n 3.27348e-19 $X=4.545 $Y=0.74 $X2=0 $Y2=0
cc_319 A1 N_A_751_74#_c_921_n 0.0193957f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_320 N_A1_c_330_n N_A_751_74#_c_921_n 0.00527124f $X=4.53 $Y=1.667 $X2=0 $Y2=0
cc_321 N_A1_M1014_g N_A_1010_74#_c_958_n 6.59741e-19 $X=4.545 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A2_c_389_n N_A3_c_442_n 0.0280268f $X=5.655 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_323 A2 A3 0.0227163f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_324 N_A2_c_387_n A3 0.00230855f $X=5.405 $Y=1.667 $X2=0 $Y2=0
cc_325 A2 N_A3_c_441_n 6.88165e-19 $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_326 N_A2_c_387_n N_A3_c_441_n 0.0111149f $X=5.405 $Y=1.667 $X2=0 $Y2=0
cc_327 N_A2_c_388_n N_A_27_392#_c_544_n 0.0129132f $X=5.205 $Y=1.885 $X2=0 $Y2=0
cc_328 A2 N_A_27_392#_c_544_n 0.0268927f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_329 N_A2_c_387_n N_A_27_392#_c_544_n 0.00611475f $X=5.405 $Y=1.667 $X2=0
+ $Y2=0
cc_330 N_A2_c_388_n N_A_27_392#_c_545_n 0.010684f $X=5.205 $Y=1.885 $X2=0 $Y2=0
cc_331 N_A2_c_389_n N_A_27_392#_c_545_n 0.0103138f $X=5.655 $Y=1.885 $X2=0 $Y2=0
cc_332 N_A2_c_389_n N_A_27_392#_c_546_n 0.0134137f $X=5.655 $Y=1.885 $X2=0 $Y2=0
cc_333 A2 N_A_27_392#_c_546_n 0.00282261f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_334 N_A2_c_387_n N_A_27_392#_c_546_n 4.5055e-19 $X=5.405 $Y=1.667 $X2=0 $Y2=0
cc_335 N_A2_c_389_n N_A_27_392#_c_547_n 6.63528e-19 $X=5.655 $Y=1.885 $X2=0
+ $Y2=0
cc_336 N_A2_c_388_n N_A_27_392#_c_552_n 5.56417e-19 $X=5.205 $Y=1.885 $X2=0
+ $Y2=0
cc_337 N_A2_c_389_n N_A_27_392#_c_552_n 5.56417e-19 $X=5.655 $Y=1.885 $X2=0
+ $Y2=0
cc_338 A2 N_A_27_392#_c_552_n 0.0276944f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_339 N_A2_c_387_n N_A_27_392#_c_552_n 0.00757755f $X=5.405 $Y=1.667 $X2=0
+ $Y2=0
cc_340 N_A2_c_388_n N_VPWR_c_676_n 0.0072484f $X=5.205 $Y=1.885 $X2=0 $Y2=0
cc_341 N_A2_c_389_n N_VPWR_c_677_n 0.00598632f $X=5.655 $Y=1.885 $X2=0 $Y2=0
cc_342 N_A2_c_388_n N_VPWR_c_686_n 0.00445602f $X=5.205 $Y=1.885 $X2=0 $Y2=0
cc_343 N_A2_c_389_n N_VPWR_c_686_n 0.00445602f $X=5.655 $Y=1.885 $X2=0 $Y2=0
cc_344 N_A2_c_388_n N_VPWR_c_672_n 0.00858665f $X=5.205 $Y=1.885 $X2=0 $Y2=0
cc_345 N_A2_c_389_n N_VPWR_c_672_n 0.00857825f $X=5.655 $Y=1.885 $X2=0 $Y2=0
cc_346 N_A2_M1011_g N_VGND_c_829_n 0.00288916f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_347 N_A2_M1026_g N_VGND_c_829_n 0.00288893f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_348 N_A2_M1011_g N_VGND_c_831_n 0.00357288f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_349 N_A2_M1026_g N_VGND_c_831_n 0.00362175f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_350 N_A2_M1011_g N_A_751_74#_c_919_n 4.10887e-19 $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_351 N_A2_M1011_g N_A_751_74#_c_920_n 0.0148139f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_352 N_A2_M1026_g N_A_751_74#_c_920_n 0.010532f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A2_M1011_g N_A_751_74#_c_922_n 4.5114e-19 $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A2_M1026_g N_A_751_74#_c_922_n 0.00682412f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A2_M1011_g N_A_1010_74#_c_960_n 0.00381522f $X=4.975 $Y=0.74 $X2=0
+ $Y2=0
cc_356 N_A2_M1026_g N_A_1010_74#_c_957_n 0.0139364f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_357 A2 N_A_1010_74#_c_957_n 0.0263457f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_358 N_A2_c_387_n N_A_1010_74#_c_957_n 0.00341628f $X=5.405 $Y=1.667 $X2=0
+ $Y2=0
cc_359 N_A2_M1011_g N_A_1010_74#_c_958_n 0.00535465f $X=4.975 $Y=0.74 $X2=0
+ $Y2=0
cc_360 A2 N_A_1010_74#_c_958_n 0.0213113f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_361 N_A2_c_387_n N_A_1010_74#_c_958_n 0.00270093f $X=5.405 $Y=1.667 $X2=0
+ $Y2=0
cc_362 N_A2_M1026_g N_A_1205_74#_c_983_n 0.00241614f $X=5.405 $Y=0.74 $X2=0
+ $Y2=0
cc_363 N_A3_c_443_n N_A4_c_500_n 0.0250804f $X=6.705 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_364 N_A3_M1018_g N_A4_M1004_g 0.0239493f $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_365 A3 A4 0.0219294f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_366 N_A3_c_441_n A4 2.27267e-19 $X=6.705 $Y=1.667 $X2=0 $Y2=0
cc_367 A3 N_A4_c_499_n 0.00350824f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_368 N_A3_c_441_n N_A4_c_499_n 0.0239528f $X=6.705 $Y=1.667 $X2=0 $Y2=0
cc_369 N_A3_c_442_n N_A_27_392#_c_545_n 6.63528e-19 $X=6.205 $Y=1.885 $X2=0
+ $Y2=0
cc_370 N_A3_c_442_n N_A_27_392#_c_546_n 0.0124513f $X=6.205 $Y=1.885 $X2=0 $Y2=0
cc_371 A3 N_A_27_392#_c_546_n 0.0289697f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_372 N_A3_c_441_n N_A_27_392#_c_546_n 4.03117e-19 $X=6.705 $Y=1.667 $X2=0
+ $Y2=0
cc_373 N_A3_c_442_n N_A_27_392#_c_547_n 0.0103043f $X=6.205 $Y=1.885 $X2=0 $Y2=0
cc_374 N_A3_c_443_n N_A_27_392#_c_547_n 0.00464047f $X=6.705 $Y=1.885 $X2=0
+ $Y2=0
cc_375 N_A3_c_443_n N_A_27_392#_c_548_n 0.0153714f $X=6.705 $Y=1.885 $X2=0 $Y2=0
cc_376 A3 N_A_27_392#_c_548_n 0.0362601f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_377 N_A3_c_441_n N_A_27_392#_c_548_n 0.00366903f $X=6.705 $Y=1.667 $X2=0
+ $Y2=0
cc_378 N_A3_c_443_n N_A_27_392#_c_550_n 5.34138e-19 $X=6.705 $Y=1.885 $X2=0
+ $Y2=0
cc_379 N_A3_c_442_n N_A_27_392#_c_553_n 5.71056e-19 $X=6.205 $Y=1.885 $X2=0
+ $Y2=0
cc_380 A3 N_A_27_392#_c_553_n 0.0277622f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_381 N_A3_c_441_n N_A_27_392#_c_553_n 0.0083547f $X=6.705 $Y=1.667 $X2=0 $Y2=0
cc_382 N_A3_c_442_n N_VPWR_c_677_n 0.00598632f $X=6.205 $Y=1.885 $X2=0 $Y2=0
cc_383 N_A3_c_442_n N_VPWR_c_678_n 5.07678e-19 $X=6.205 $Y=1.885 $X2=0 $Y2=0
cc_384 N_A3_c_443_n N_VPWR_c_678_n 0.0108529f $X=6.705 $Y=1.885 $X2=0 $Y2=0
cc_385 N_A3_c_442_n N_VPWR_c_687_n 0.00445602f $X=6.205 $Y=1.885 $X2=0 $Y2=0
cc_386 N_A3_c_443_n N_VPWR_c_687_n 0.00413917f $X=6.705 $Y=1.885 $X2=0 $Y2=0
cc_387 N_A3_c_442_n N_VPWR_c_672_n 0.00858286f $X=6.205 $Y=1.885 $X2=0 $Y2=0
cc_388 N_A3_c_443_n N_VPWR_c_672_n 0.00818187f $X=6.705 $Y=1.885 $X2=0 $Y2=0
cc_389 N_A3_M1018_g N_VGND_c_826_n 3.70941e-19 $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_390 N_A3_M1007_g N_VGND_c_829_n 0.00278247f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A3_M1018_g N_VGND_c_829_n 0.00278247f $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A3_M1007_g N_VGND_c_831_n 0.00358425f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_393 N_A3_M1018_g N_VGND_c_831_n 0.00353524f $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_394 N_A3_M1007_g N_A_751_74#_c_922_n 6.27938e-19 $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_395 N_A3_M1007_g N_A_1010_74#_c_957_n 0.0158982f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_396 N_A3_M1018_g N_A_1010_74#_c_957_n 0.00140095f $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_397 A3 N_A_1010_74#_c_957_n 0.0616708f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_398 N_A3_c_441_n N_A_1010_74#_c_957_n 0.0072954f $X=6.705 $Y=1.667 $X2=0
+ $Y2=0
cc_399 N_A3_M1007_g N_A_1205_74#_c_981_n 0.00684765f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_400 N_A3_M1018_g N_A_1205_74#_c_981_n 5.91819e-19 $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A3_M1007_g N_A_1205_74#_c_982_n 0.0100245f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_402 N_A3_M1018_g N_A_1205_74#_c_982_n 0.0116238f $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_403 N_A3_M1007_g N_A_1205_74#_c_983_n 0.00281658f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_404 N_A3_M1007_g N_A_1205_74#_c_993_n 6.44259e-19 $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_405 N_A3_M1018_g N_A_1205_74#_c_993_n 0.00880957f $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A3_M1018_g N_A_1205_74#_c_985_n 0.0040946f $X=6.81 $Y=0.74 $X2=0 $Y2=0
cc_407 A3 N_A_1205_74#_c_985_n 0.0188033f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_408 N_A4_c_500_n N_A_27_392#_c_548_n 0.0141516f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_409 N_A4_c_499_n N_A_27_392#_c_548_n 4.92109e-19 $X=7.655 $Y=1.667 $X2=0
+ $Y2=0
cc_410 N_A4_c_500_n N_A_27_392#_c_549_n 8.00885e-19 $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_411 N_A4_c_501_n N_A_27_392#_c_549_n 0.00216588f $X=7.655 $Y=1.885 $X2=0
+ $Y2=0
cc_412 A4 N_A_27_392#_c_549_n 0.0227022f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_413 N_A4_c_499_n N_A_27_392#_c_549_n 0.00821828f $X=7.655 $Y=1.667 $X2=0
+ $Y2=0
cc_414 N_A4_c_500_n N_A_27_392#_c_550_n 0.010218f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_415 N_A4_c_501_n N_A_27_392#_c_550_n 0.00960826f $X=7.655 $Y=1.885 $X2=0
+ $Y2=0
cc_416 N_A4_c_500_n N_VPWR_c_678_n 0.0068696f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_417 N_A4_c_501_n N_VPWR_c_680_n 0.008504f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_418 A4 N_VPWR_c_680_n 0.0211423f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_419 N_A4_c_500_n N_VPWR_c_688_n 0.00445602f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_420 N_A4_c_501_n N_VPWR_c_688_n 0.00445602f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_421 N_A4_c_500_n N_VPWR_c_672_n 0.00857432f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_422 N_A4_c_501_n N_VPWR_c_672_n 0.00861084f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_423 N_A4_M1004_g N_VGND_c_826_n 0.00974368f $X=7.24 $Y=0.74 $X2=0 $Y2=0
cc_424 N_A4_M1015_g N_VGND_c_826_n 0.0133215f $X=7.67 $Y=0.74 $X2=0 $Y2=0
cc_425 N_A4_M1004_g N_VGND_c_829_n 0.00383152f $X=7.24 $Y=0.74 $X2=0 $Y2=0
cc_426 N_A4_M1015_g N_VGND_c_830_n 0.00383152f $X=7.67 $Y=0.74 $X2=0 $Y2=0
cc_427 N_A4_M1004_g N_VGND_c_831_n 0.00757637f $X=7.24 $Y=0.74 $X2=0 $Y2=0
cc_428 N_A4_M1015_g N_VGND_c_831_n 0.0076118f $X=7.67 $Y=0.74 $X2=0 $Y2=0
cc_429 N_A4_M1004_g N_A_1205_74#_c_982_n 9.48753e-19 $X=7.24 $Y=0.74 $X2=0 $Y2=0
cc_430 N_A4_M1004_g N_A_1205_74#_c_984_n 0.0163723f $X=7.24 $Y=0.74 $X2=0 $Y2=0
cc_431 N_A4_M1015_g N_A_1205_74#_c_984_n 0.0157274f $X=7.67 $Y=0.74 $X2=0 $Y2=0
cc_432 A4 N_A_1205_74#_c_984_n 0.0562102f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_433 N_A4_c_499_n N_A_1205_74#_c_984_n 0.00376693f $X=7.655 $Y=1.667 $X2=0
+ $Y2=0
cc_434 N_A4_M1015_g N_A_1205_74#_c_986_n 0.00160885f $X=7.67 $Y=0.74 $X2=0 $Y2=0
cc_435 N_A_27_392#_c_542_n N_VPWR_M1000_d 0.00777378f $X=4.045 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_436 N_A_27_392#_c_542_n N_VPWR_M1001_d 0.00379433f $X=4.045 $Y=2.375 $X2=0
+ $Y2=0
cc_437 N_A_27_392#_c_542_n N_VPWR_M1027_d 0.00761902f $X=4.045 $Y=2.375 $X2=0
+ $Y2=0
cc_438 N_A_27_392#_c_544_n N_VPWR_M1008_d 0.00582112f $X=5.265 $Y=2.035 $X2=0
+ $Y2=0
cc_439 N_A_27_392#_c_546_n N_VPWR_M1025_s 0.00339226f $X=6.265 $Y=2.035 $X2=0
+ $Y2=0
cc_440 N_A_27_392#_c_548_n N_VPWR_M1021_d 0.00250873f $X=7.265 $Y=2.035 $X2=0
+ $Y2=0
cc_441 N_A_27_392#_c_538_n N_VPWR_c_673_n 0.0121617f $X=1.065 $Y=2.99 $X2=0
+ $Y2=0
cc_442 N_A_27_392#_c_541_n N_VPWR_c_673_n 0.0185064f $X=1.23 $Y=2.815 $X2=0
+ $Y2=0
cc_443 N_A_27_392#_c_542_n N_VPWR_c_673_n 0.0219924f $X=4.045 $Y=2.375 $X2=0
+ $Y2=0
cc_444 N_A_27_392#_c_542_n N_VPWR_c_674_n 0.0171814f $X=4.045 $Y=2.375 $X2=0
+ $Y2=0
cc_445 N_A_27_392#_c_542_n N_VPWR_c_675_n 0.0201047f $X=4.045 $Y=2.375 $X2=0
+ $Y2=0
cc_446 N_A_27_392#_c_551_n N_VPWR_c_675_n 0.0100206f $X=4.21 $Y=2.455 $X2=0
+ $Y2=0
cc_447 N_A_27_392#_c_544_n N_VPWR_c_676_n 0.0334384f $X=5.265 $Y=2.035 $X2=0
+ $Y2=0
cc_448 N_A_27_392#_c_545_n N_VPWR_c_676_n 0.0267216f $X=5.43 $Y=2.815 $X2=0
+ $Y2=0
cc_449 N_A_27_392#_c_551_n N_VPWR_c_676_n 0.0158658f $X=4.21 $Y=2.455 $X2=0
+ $Y2=0
cc_450 N_A_27_392#_c_545_n N_VPWR_c_677_n 0.0266809f $X=5.43 $Y=2.815 $X2=0
+ $Y2=0
cc_451 N_A_27_392#_c_546_n N_VPWR_c_677_n 0.0232685f $X=6.265 $Y=2.035 $X2=0
+ $Y2=0
cc_452 N_A_27_392#_c_547_n N_VPWR_c_677_n 0.0266809f $X=6.43 $Y=2.815 $X2=0
+ $Y2=0
cc_453 N_A_27_392#_c_547_n N_VPWR_c_678_n 0.0266809f $X=6.43 $Y=2.815 $X2=0
+ $Y2=0
cc_454 N_A_27_392#_c_548_n N_VPWR_c_678_n 0.0202249f $X=7.265 $Y=2.035 $X2=0
+ $Y2=0
cc_455 N_A_27_392#_c_550_n N_VPWR_c_678_n 0.0266809f $X=7.43 $Y=2.815 $X2=0
+ $Y2=0
cc_456 N_A_27_392#_c_549_n N_VPWR_c_680_n 0.0121172f $X=7.43 $Y=2.12 $X2=0 $Y2=0
cc_457 N_A_27_392#_c_550_n N_VPWR_c_680_n 0.0576605f $X=7.43 $Y=2.815 $X2=0
+ $Y2=0
cc_458 N_A_27_392#_c_551_n N_VPWR_c_681_n 0.0146357f $X=4.21 $Y=2.455 $X2=0
+ $Y2=0
cc_459 N_A_27_392#_c_538_n N_VPWR_c_683_n 0.0627048f $X=1.065 $Y=2.99 $X2=0
+ $Y2=0
cc_460 N_A_27_392#_c_539_n N_VPWR_c_683_n 0.0236039f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_461 N_A_27_392#_c_545_n N_VPWR_c_686_n 0.014552f $X=5.43 $Y=2.815 $X2=0 $Y2=0
cc_462 N_A_27_392#_c_547_n N_VPWR_c_687_n 0.0145938f $X=6.43 $Y=2.815 $X2=0
+ $Y2=0
cc_463 N_A_27_392#_c_550_n N_VPWR_c_688_n 0.014552f $X=7.43 $Y=2.815 $X2=0 $Y2=0
cc_464 N_A_27_392#_c_538_n N_VPWR_c_672_n 0.0348361f $X=1.065 $Y=2.99 $X2=0
+ $Y2=0
cc_465 N_A_27_392#_c_539_n N_VPWR_c_672_n 0.012761f $X=0.445 $Y=2.99 $X2=0 $Y2=0
cc_466 N_A_27_392#_c_545_n N_VPWR_c_672_n 0.0119791f $X=5.43 $Y=2.815 $X2=0
+ $Y2=0
cc_467 N_A_27_392#_c_547_n N_VPWR_c_672_n 0.0120466f $X=6.43 $Y=2.815 $X2=0
+ $Y2=0
cc_468 N_A_27_392#_c_550_n N_VPWR_c_672_n 0.0119791f $X=7.43 $Y=2.815 $X2=0
+ $Y2=0
cc_469 N_A_27_392#_c_551_n N_VPWR_c_672_n 0.0121141f $X=4.21 $Y=2.455 $X2=0
+ $Y2=0
cc_470 N_A_27_392#_c_542_n N_X_M1000_s 0.00891825f $X=4.045 $Y=2.375 $X2=0 $Y2=0
cc_471 N_A_27_392#_c_542_n N_X_M1003_s 0.00891405f $X=4.045 $Y=2.375 $X2=0 $Y2=0
cc_472 N_A_27_392#_c_542_n N_X_c_790_n 0.0255897f $X=4.045 $Y=2.375 $X2=0 $Y2=0
cc_473 N_A_27_392#_c_542_n N_X_c_805_n 0.0427079f $X=4.045 $Y=2.375 $X2=0 $Y2=0
cc_474 N_A_27_392#_c_546_n N_A_1010_74#_c_957_n 0.00685685f $X=6.265 $Y=2.035
+ $X2=0 $Y2=0
cc_475 N_A_27_392#_c_548_n N_A_1205_74#_c_984_n 0.00357224f $X=7.265 $Y=2.035
+ $X2=0 $Y2=0
cc_476 N_A_27_392#_c_549_n N_A_1205_74#_c_984_n 0.00167234f $X=7.43 $Y=2.12
+ $X2=0 $Y2=0
cc_477 N_A_27_392#_c_548_n N_A_1205_74#_c_985_n 0.00113065f $X=7.265 $Y=2.035
+ $X2=0 $Y2=0
cc_478 N_VPWR_M1001_d N_X_c_805_n 0.00206339f $X=2.54 $Y=1.84 $X2=0 $Y2=0
cc_479 N_VPWR_c_680_n N_A_1205_74#_c_984_n 3.21545e-19 $X=7.88 $Y=2.115 $X2=0
+ $Y2=0
cc_480 N_X_c_783_n N_VGND_M1009_d 0.00664343f $X=2.555 $Y=1.085 $X2=0 $Y2=0
cc_481 N_X_c_794_n N_VGND_M1023_d 0.00744145f $X=2.93 $Y=1.17 $X2=0 $Y2=0
cc_482 X N_VGND_M1023_d 0.00266152f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_483 N_X_c_794_n N_A_751_74#_c_921_n 0.00599151f $X=2.93 $Y=1.17 $X2=0 $Y2=0
cc_484 N_VGND_c_831_n N_A_751_74#_c_917_n 0.00734594f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_485 N_VGND_c_829_n N_A_751_74#_c_918_n 0.00824596f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_486 N_VGND_c_831_n N_A_751_74#_c_918_n 0.00635316f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_c_829_n N_A_751_74#_c_920_n 0.0267924f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_488 N_VGND_c_831_n N_A_751_74#_c_920_n 0.0208291f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_489 N_VGND_c_829_n N_A_751_74#_c_922_n 0.0158045f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_490 N_VGND_c_831_n N_A_751_74#_c_922_n 0.01217f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_491 N_VGND_c_826_n N_A_1205_74#_c_982_n 0.0112234f $X=7.455 $Y=0.495 $X2=0
+ $Y2=0
cc_492 N_VGND_c_829_n N_A_1205_74#_c_982_n 0.0511953f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_493 N_VGND_c_831_n N_A_1205_74#_c_982_n 0.0283873f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_494 N_VGND_c_829_n N_A_1205_74#_c_983_n 0.0235818f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_495 N_VGND_c_831_n N_A_1205_74#_c_983_n 0.0127177f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_496 N_VGND_c_826_n N_A_1205_74#_c_984_n 0.0216087f $X=7.455 $Y=0.495 $X2=0
+ $Y2=0
cc_497 N_VGND_c_826_n N_A_1205_74#_c_986_n 0.0229007f $X=7.455 $Y=0.495 $X2=0
+ $Y2=0
cc_498 N_VGND_c_830_n N_A_1205_74#_c_986_n 0.0115122f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_499 N_VGND_c_831_n N_A_1205_74#_c_986_n 0.0095288f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_500 N_A_751_74#_c_920_n N_A_1010_74#_M1011_s 0.00178994f $X=5.455 $Y=0.465
+ $X2=-0.19 $Y2=-0.245
cc_501 N_A_751_74#_c_920_n N_A_1010_74#_c_960_n 0.0149186f $X=5.455 $Y=0.465
+ $X2=0 $Y2=0
cc_502 N_A_751_74#_c_920_n N_A_1010_74#_c_957_n 0.004342f $X=5.455 $Y=0.465
+ $X2=0 $Y2=0
cc_503 N_A_751_74#_c_922_n N_A_1010_74#_c_957_n 0.0242226f $X=5.62 $Y=0.515
+ $X2=0 $Y2=0
cc_504 N_A_751_74#_c_919_n N_A_1010_74#_c_958_n 0.00336899f $X=4.76 $Y=0.77
+ $X2=0 $Y2=0
cc_505 N_A_751_74#_c_922_n N_A_1205_74#_c_981_n 0.0370692f $X=5.62 $Y=0.515
+ $X2=0 $Y2=0
cc_506 N_A_751_74#_c_922_n N_A_1205_74#_c_983_n 0.00753743f $X=5.62 $Y=0.515
+ $X2=0 $Y2=0
cc_507 N_A_1010_74#_c_957_n N_A_1205_74#_c_981_n 0.0244212f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_508 N_A_1010_74#_M1007_s N_A_1205_74#_c_982_n 0.00176461f $X=6.455 $Y=0.37
+ $X2=0 $Y2=0
cc_509 N_A_1010_74#_c_979_p N_A_1205_74#_c_982_n 0.0126419f $X=6.595 $Y=0.785
+ $X2=0 $Y2=0
cc_510 N_A_1010_74#_c_957_n N_A_1205_74#_c_985_n 0.0144643f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
