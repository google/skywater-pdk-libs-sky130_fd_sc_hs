* File: sky130_fd_sc_hs__diode_2.spice
* Created: Thu Aug 27 20:40:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__diode_2.pex.spice"
.subckt sky130_fd_sc_hs__diode_2  VNB VPB DIODE VGND VPWR
* 
* DIODE	DIODE
* VPB	VPB
* VNB	VNB
D0_noxref VNB N_DIODE_D0_noxref_neg NDIODE  AREA=0.6417 PJ=3.24 M=1
+ AHFTEMPPERIM=3.24
DX1_noxref VNB VPB NWDIODE A=2.4924 P=6.4
*
.include "sky130_fd_sc_hs__diode_2.pxi.spice"
*
.ends
*
*
