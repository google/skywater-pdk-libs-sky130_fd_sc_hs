* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__or2b_1 A B_N VGND VNB VPB VPWR X
M1000 a_264_368# a_27_112# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=7.357e+11p ps=5.01e+06u
M1001 VGND A a_264_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND B_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=3.685e+11p ps=2.44e+06u
M1003 X a_264_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=7.662e+11p ps=5.48e+06u
M1004 a_353_368# a_27_112# a_264_368# VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=2.95e+11p ps=2.59e+06u
M1005 VPWR B_N a_27_112# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1006 VPWR A a_353_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_264_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends
