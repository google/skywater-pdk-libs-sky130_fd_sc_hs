* File: sky130_fd_sc_hs__a32o_4.pex.spice
* Created: Thu Aug 27 20:30:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A32O_4%A_83_283# 1 2 3 4 13 15 16 18 19 21 22 24 25
+ 27 30 32 34 37 39 48 49 50 53 56 59 60 62 67 69 81
c177 69 0 1.2831e-19 $X=5.965 $Y=1.1
c178 67 0 7.34128e-20 $X=4.19 $Y=2.115
c179 60 0 7.32746e-20 $X=4.055 $Y=1.195
c180 59 0 1.79774e-20 $X=5.8 $Y=1.195
r181 75 76 1.83038 $w=3.95e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.515
+ $X2=0.955 $Y2=1.515
r182 74 75 53.081 $w=3.95e-07 $l=4.35e-07 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.94 $Y2=1.515
r183 73 74 1.22025 $w=3.95e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.505 $Y2=1.515
r184 69 71 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.965 $Y=1.1
+ $X2=5.965 $Y2=1.195
r185 64 65 26.5367 $w=1.77e-07 $l=3.85e-07 $layer=LI1_cond $X=3.585 $Y=1.187
+ $X2=3.97 $Y2=1.187
r186 60 65 5.85876 $w=1.77e-07 $l=8.89101e-08 $layer=LI1_cond $X=4.055 $Y=1.195
+ $X2=3.97 $Y2=1.187
r187 59 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.8 $Y=1.195
+ $X2=5.965 $Y2=1.195
r188 59 60 113.845 $w=1.68e-07 $l=1.745e-06 $layer=LI1_cond $X=5.8 $Y=1.195
+ $X2=4.055 $Y2=1.195
r189 56 67 3.70735 $w=2.5e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.97 $Y=1.95
+ $X2=4.12 $Y2=2.035
r190 55 65 0.961343 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=3.97 $Y=1.28
+ $X2=3.97 $Y2=1.187
r191 55 56 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.97 $Y=1.28
+ $X2=3.97 $Y2=1.95
r192 54 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=2.035
+ $X2=3.19 $Y2=2.035
r193 53 67 2.76166 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.885 $Y=2.035
+ $X2=4.12 $Y2=2.035
r194 53 54 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.885 $Y=2.035
+ $X2=3.355 $Y2=2.035
r195 49 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=2.035
+ $X2=3.19 $Y2=2.035
r196 49 50 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.025 $Y=2.035
+ $X2=2.185 $Y2=2.035
r197 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.1 $Y=1.95
+ $X2=2.185 $Y2=2.035
r198 47 48 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.1 $Y=1.68 $X2=2.1
+ $Y2=1.95
r199 46 81 9.1519 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.515
+ $X2=1.905 $Y2=1.515
r200 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.515 $X2=1.83 $Y2=1.515
r201 42 78 37.2177 $w=3.95e-07 $l=3.05e-07 $layer=POLY_cond $X=1.15 $Y=1.515
+ $X2=1.455 $Y2=1.515
r202 42 76 23.7949 $w=3.95e-07 $l=1.95e-07 $layer=POLY_cond $X=1.15 $Y=1.515
+ $X2=0.955 $Y2=1.515
r203 41 45 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.15 $Y=1.515
+ $X2=1.83 $Y2=1.515
r204 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.515 $X2=1.15 $Y2=1.515
r205 39 47 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.015 $Y=1.515
+ $X2=2.1 $Y2=1.68
r206 39 45 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.015 $Y=1.515
+ $X2=1.83 $Y2=1.515
r207 35 81 5.49114 $w=3.95e-07 $l=4.5e-08 $layer=POLY_cond $X=1.95 $Y=1.515
+ $X2=1.905 $Y2=1.515
r208 35 37 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.95 $Y=1.35
+ $X2=1.95 $Y2=0.82
r209 32 81 25.5547 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=1.515
r210 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=2.4
r211 28 46 37.8278 $w=3.95e-07 $l=3.1e-07 $layer=POLY_cond $X=1.52 $Y=1.515
+ $X2=1.83 $Y2=1.515
r212 28 78 7.93165 $w=3.95e-07 $l=6.5e-08 $layer=POLY_cond $X=1.52 $Y=1.515
+ $X2=1.455 $Y2=1.515
r213 28 30 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.52 $Y=1.35
+ $X2=1.52 $Y2=0.82
r214 25 78 25.5547 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.515
r215 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r216 22 76 25.5547 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.515
r217 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r218 19 75 25.5547 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.94 $Y=1.265
+ $X2=0.94 $Y2=1.515
r219 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.94 $Y=1.265
+ $X2=0.94 $Y2=0.82
r220 16 74 25.5547 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.515
r221 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r222 13 73 25.5547 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.495 $Y=1.265
+ $X2=0.495 $Y2=1.515
r223 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.265
+ $X2=0.495 $Y2=0.82
r224 4 67 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=1.96 $X2=4.19 $Y2=2.115
r225 3 62 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=2.99
+ $Y=1.96 $X2=3.19 $Y2=2.115
r226 2 69 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.825
+ $Y=0.61 $X2=5.965 $Y2=1.1
r227 1 64 182 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.55 $X2=3.585 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%B2 3 5 7 8 10 11 13 14 17 19 20 24 28 29 30
+ 36 44 46
c107 44 0 6.39601e-20 $X=4.415 $Y=0.42
c108 30 0 1.33336e-19 $X=4.25 $Y=0.34
c109 19 0 1.0936e-19 $X=4.81 $Y=1.08
c110 11 0 7.39242e-20 $X=4.415 $Y=1.885
c111 8 0 7.32746e-20 $X=4.23 $Y=0.585
r112 36 46 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=1.615
+ $X2=2.67 $Y2=1.45
r113 36 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.615 $X2=2.67 $Y2=1.615
r114 34 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=0.42
+ $X2=4.415 $Y2=0.42
r115 34 41 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.25 $Y=0.42 $X2=4.23
+ $Y2=0.42
r116 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.25
+ $Y=0.42 $X2=4.25 $Y2=0.42
r117 30 33 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.25 $Y=0.34 $X2=4.25
+ $Y2=0.42
r118 28 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=0.34
+ $X2=4.25 $Y2=0.34
r119 28 29 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=4.085 $Y=0.34
+ $X2=2.74 $Y2=0.34
r120 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.655 $Y=0.425
+ $X2=2.74 $Y2=0.34
r121 26 46 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.655 $Y=0.425
+ $X2=2.655 $Y2=1.45
r122 22 24 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=4.705 $Y=1.155
+ $X2=4.81 $Y2=1.155
r123 20 21 86.8199 $w=1.61e-07 $l=2.9e-07 $layer=POLY_cond $X=4.415 $Y=1.795
+ $X2=4.705 $Y2=1.795
r124 19 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.81 $Y=1.08
+ $X2=4.81 $Y2=1.155
r125 18 19 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.81 $Y=0.585
+ $X2=4.81 $Y2=1.08
r126 17 21 4.52116 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.705 $Y=1.705
+ $X2=4.705 $Y2=1.795
r127 16 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=1.23
+ $X2=4.705 $Y2=1.155
r128 16 17 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.705 $Y=1.23
+ $X2=4.705 $Y2=1.705
r129 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.735 $Y=0.51
+ $X2=4.81 $Y2=0.585
r130 14 44 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.735 $Y=0.51
+ $X2=4.415 $Y2=0.51
r131 11 20 4.52116 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.415 $Y=1.885
+ $X2=4.415 $Y2=1.795
r132 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.415 $Y=1.885
+ $X2=4.415 $Y2=2.46
r133 8 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=0.585
+ $X2=4.23 $Y2=0.42
r134 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.23 $Y=0.585
+ $X2=4.23 $Y2=1.015
r135 5 39 52.0344 $w=4.22e-07 $l=3.40734e-07 $layer=POLY_cond $X=2.915 $Y=1.885
+ $X2=2.755 $Y2=1.615
r136 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.915 $Y=1.885
+ $X2=2.915 $Y2=2.46
r137 1 39 40.0415 $w=4.22e-07 $l=2.11069e-07 $layer=POLY_cond $X=2.86 $Y=1.45
+ $X2=2.755 $Y2=1.615
r138 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.86 $Y=1.45 $X2=2.86
+ $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%B1 3 5 7 8 10 11 13 14 15 23
c56 23 0 8.37829e-20 $X=3.8 $Y=1.667
c57 8 0 1.33336e-19 $X=3.8 $Y=1.45
r58 21 23 43.8182 $w=3.41e-07 $l=3.1e-07 $layer=POLY_cond $X=3.49 $Y=1.667
+ $X2=3.8 $Y2=1.667
r59 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.615 $X2=3.49 $Y2=1.615
r60 19 21 10.6012 $w=3.41e-07 $l=7.5e-08 $layer=POLY_cond $X=3.415 $Y=1.667
+ $X2=3.49 $Y2=1.667
r61 15 22 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.6 $Y=1.615
+ $X2=3.49 $Y2=1.615
r62 14 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.615
+ $X2=3.49 $Y2=1.615
r63 11 23 16.2551 $w=3.41e-07 $l=2.69433e-07 $layer=POLY_cond $X=3.915 $Y=1.885
+ $X2=3.8 $Y2=1.667
r64 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.915 $Y=1.885
+ $X2=3.915 $Y2=2.46
r65 8 23 22.0049 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=3.8 $Y=1.45 $X2=3.8
+ $Y2=1.667
r66 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.8 $Y=1.45 $X2=3.8
+ $Y2=1.015
r67 5 19 22.0049 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=3.415 $Y=1.885
+ $X2=3.415 $Y2=1.667
r68 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.415 $Y=1.885
+ $X2=3.415 $Y2=2.46
r69 1 19 17.6686 $w=3.41e-07 $l=2.72422e-07 $layer=POLY_cond $X=3.29 $Y=1.45
+ $X2=3.415 $Y2=1.667
r70 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.29 $Y=1.45 $X2=3.29
+ $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%A2 1 3 6 10 12 14 15 16 17 18 20 21 28 31
c105 28 0 6.33061e-20 $X=6.66 $Y=1.605
c106 21 0 8.37829e-20 $X=5.18 $Y=1.63
c107 18 0 7.39242e-20 $X=5.35 $Y=2.035
c108 10 0 3.2498e-19 $X=6.69 $Y=0.93
c109 6 0 1.13206e-20 $X=5.32 $Y=0.93
c110 1 0 7.34128e-20 $X=5.11 $Y=1.885
r111 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.605 $X2=6.66 $Y2=1.605
r112 25 28 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.51 $Y=1.605
+ $X2=6.66 $Y2=1.605
r113 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.185
+ $Y=1.635 $X2=5.185 $Y2=1.635
r114 21 31 5.3375 $w=3.2e-07 $l=1.4e-07 $layer=LI1_cond $X=5.18 $Y=1.63 $X2=5.04
+ $Y2=1.63
r115 21 23 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=1.63
+ $X2=5.265 $Y2=1.63
r116 19 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.51 $Y=1.77
+ $X2=6.51 $Y2=1.605
r117 19 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.51 $Y=1.77
+ $X2=6.51 $Y2=1.95
r118 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=6.51 $Y2=1.95
r119 17 18 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=5.35 $Y2=2.035
r120 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.265 $Y=1.95
+ $X2=5.35 $Y2=2.035
r121 15 23 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.265 $Y=1.79
+ $X2=5.265 $Y2=1.63
r122 15 16 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.265 $Y=1.79
+ $X2=5.265 $Y2=1.95
r123 12 29 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=6.705 $Y=1.885
+ $X2=6.66 $Y2=1.605
r124 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.705 $Y=1.885
+ $X2=6.705 $Y2=2.46
r125 8 29 38.6072 $w=2.91e-07 $l=1.79374e-07 $layer=POLY_cond $X=6.69 $Y=1.44
+ $X2=6.66 $Y2=1.605
r126 8 10 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.69 $Y=1.44
+ $X2=6.69 $Y2=0.93
r127 4 24 38.6365 $w=3.35e-07 $l=2.14173e-07 $layer=POLY_cond $X=5.32 $Y=1.47
+ $X2=5.207 $Y2=1.635
r128 4 6 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.32 $Y=1.47 $X2=5.32
+ $Y2=0.93
r129 1 24 50.8664 $w=3.35e-07 $l=2.94534e-07 $layer=POLY_cond $X=5.11 $Y=1.885
+ $X2=5.207 $Y2=1.635
r130 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.11 $Y=1.885
+ $X2=5.11 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%A1 1 3 6 10 12 14 15 22
c55 12 0 1.12995e-19 $X=6.195 $Y=1.885
c56 10 0 1.83396e-19 $X=6.18 $Y=0.93
c57 6 0 2.77406e-20 $X=5.75 $Y=0.93
r58 22 23 1.8634 $w=3.88e-07 $l=1.5e-08 $layer=POLY_cond $X=6.18 $Y=1.667
+ $X2=6.195 $Y2=1.667
r59 20 22 47.2062 $w=3.88e-07 $l=3.8e-07 $layer=POLY_cond $X=5.8 $Y=1.667
+ $X2=6.18 $Y2=1.667
r60 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.8
+ $Y=1.615 $X2=5.8 $Y2=1.615
r61 18 20 6.21134 $w=3.88e-07 $l=5e-08 $layer=POLY_cond $X=5.75 $Y=1.667 $X2=5.8
+ $Y2=1.667
r62 17 18 3.10567 $w=3.88e-07 $l=2.5e-08 $layer=POLY_cond $X=5.725 $Y=1.667
+ $X2=5.75 $Y2=1.667
r63 15 21 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6 $Y=1.615 $X2=5.8
+ $Y2=1.615
r64 12 23 25.1189 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.195 $Y=1.885
+ $X2=6.195 $Y2=1.667
r65 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.195 $Y=1.885
+ $X2=6.195 $Y2=2.46
r66 8 22 25.1189 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.18 $Y=1.45
+ $X2=6.18 $Y2=1.667
r67 8 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.18 $Y=1.45 $X2=6.18
+ $Y2=0.93
r68 4 18 25.1189 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.75 $Y=1.45
+ $X2=5.75 $Y2=1.667
r69 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.75 $Y=1.45 $X2=5.75
+ $Y2=0.93
r70 1 17 25.1189 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.725 $Y=1.885
+ $X2=5.725 $Y2=1.667
r71 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.725 $Y=1.885
+ $X2=5.725 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%A3 3 5 7 8 10 13 15 16 24
c52 3 0 6.33061e-20 $X=7.14 $Y=0.93
r53 24 25 1.26842 $w=3.8e-07 $l=1e-08 $layer=POLY_cond $X=7.655 $Y=1.667
+ $X2=7.665 $Y2=1.667
r54 22 24 0.634211 $w=3.8e-07 $l=5e-09 $layer=POLY_cond $X=7.65 $Y=1.667
+ $X2=7.655 $Y2=1.667
r55 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.65
+ $Y=1.615 $X2=7.65 $Y2=1.615
r56 20 22 62.7868 $w=3.8e-07 $l=4.95e-07 $layer=POLY_cond $X=7.155 $Y=1.667
+ $X2=7.65 $Y2=1.667
r57 19 20 1.90263 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=7.14 $Y=1.667
+ $X2=7.155 $Y2=1.667
r58 16 23 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.92 $Y=1.615
+ $X2=7.65 $Y2=1.615
r59 15 23 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.44 $Y=1.615
+ $X2=7.65 $Y2=1.615
r60 11 25 24.6126 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=7.665 $Y=1.45
+ $X2=7.665 $Y2=1.667
r61 11 13 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.665 $Y=1.45
+ $X2=7.665 $Y2=0.93
r62 8 24 24.6126 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.655 $Y=1.885
+ $X2=7.655 $Y2=1.667
r63 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.655 $Y=1.885
+ $X2=7.655 $Y2=2.46
r64 5 20 24.6126 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.155 $Y=1.885
+ $X2=7.155 $Y2=1.667
r65 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.155 $Y=1.885
+ $X2=7.155 $Y2=2.46
r66 1 19 24.6126 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=7.14 $Y=1.45
+ $X2=7.14 $Y2=1.667
r67 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.14 $Y=1.45 $X2=7.14
+ $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 39 43 45 47
+ 52 57 65 70 77 78 84 87 90 93 96
r111 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r113 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r114 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r116 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r117 78 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r119 75 96 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.405 $Y2=3.33
r120 75 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 74 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 74 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 71 93 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.645 $Y=3.33
+ $X2=6.465 $Y2=3.33
r125 71 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.645 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 70 96 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.405 $Y2=3.33
r127 70 73 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=6.96 $Y2=3.33
r128 69 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r129 69 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r130 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r131 66 90 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.615 $Y=3.33
+ $X2=5.412 $Y2=3.33
r132 66 68 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.615 $Y=3.33
+ $X2=6 $Y2=3.33
r133 65 93 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.285 $Y=3.33
+ $X2=6.465 $Y2=3.33
r134 65 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.285 $Y=3.33
+ $X2=6 $Y2=3.33
r135 64 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r136 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r137 61 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 60 63 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=5.04 $Y2=3.33
r139 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r140 58 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.13 $Y2=3.33
r141 58 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r142 57 90 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.412 $Y2=3.33
r143 57 63 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 56 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r145 56 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r146 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r147 53 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r148 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r149 52 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.13 $Y2=3.33
r150 52 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.68 $Y2=3.33
r151 51 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r152 51 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r153 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 48 81 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r155 48 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r156 47 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r157 47 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r158 45 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r159 45 61 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r160 41 96 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=3.245
+ $X2=7.405 $Y2=3.33
r161 41 43 32.5154 $w=2.78e-07 $l=7.9e-07 $layer=LI1_cond $X=7.405 $Y=3.245
+ $X2=7.405 $Y2=2.455
r162 37 93 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.465 $Y=3.245
+ $X2=6.465 $Y2=3.33
r163 37 39 14.4055 $w=3.58e-07 $l=4.5e-07 $layer=LI1_cond $X=6.465 $Y=3.245
+ $X2=6.465 $Y2=2.795
r164 33 90 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.412 $Y=3.245
+ $X2=5.412 $Y2=3.33
r165 33 35 13.9431 $w=4.03e-07 $l=4.9e-07 $layer=LI1_cond $X=5.412 $Y=3.245
+ $X2=5.412 $Y2=2.755
r166 29 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=3.33
r167 29 31 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=2.405
r168 25 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r169 25 27 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.295
r170 21 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r171 19 81 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r172 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r173 6 43 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=7.23
+ $Y=1.96 $X2=7.38 $Y2=2.455
r174 5 39 600 $w=1.7e-07 $l=9.27389e-07 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.96 $X2=6.465 $Y2=2.795
r175 4 35 600 $w=1.7e-07 $l=8.91628e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.96 $X2=5.39 $Y2=2.755
r176 3 31 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=1.98
+ $Y=1.84 $X2=2.13 $Y2=2.405
r177 2 27 300 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.295
r178 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r179 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%X 1 2 3 4 13 14 15 16 18 21 25 27 29 31 33 37
+ 42 44 47
c70 47 0 1.55137e-19 $X=0.24 $Y=1.295
c71 13 0 1.58808e-19 $X=0.615 $Y=1.055
r72 40 47 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.24 $Y=1.48
+ $X2=0.24 $Y2=1.295
r73 39 47 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.18
+ $X2=0.24 $Y2=1.295
r74 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.735 $Y=0.93
+ $X2=1.735 $Y2=0.595
r75 31 46 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=2.02
+ $X2=1.655 $Y2=1.935
r76 31 33 33.5443 $w=2.78e-07 $l=8.15e-07 $layer=LI1_cond $X=1.655 $Y=2.02
+ $X2=1.655 $Y2=2.835
r77 30 44 4.36636 $w=2.5e-07 $l=1.03e-07 $layer=LI1_cond $X=0.82 $Y=1.055
+ $X2=0.717 $Y2=1.055
r78 29 35 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=1.57 $Y=1.055
+ $X2=1.735 $Y2=0.93
r79 29 30 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=1.57 $Y=1.055
+ $X2=0.82 $Y2=1.055
r80 28 42 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=1.935
+ $X2=0.69 $Y2=1.935
r81 27 46 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.515 $Y=1.935
+ $X2=1.655 $Y2=1.935
r82 27 28 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.515 $Y=1.935
+ $X2=0.815 $Y2=1.935
r83 23 44 2.066 $w=2.05e-07 $l=1.25e-07 $layer=LI1_cond $X=0.717 $Y=0.93
+ $X2=0.717 $Y2=1.055
r84 23 25 19.2062 $w=2.03e-07 $l=3.55e-07 $layer=LI1_cond $X=0.717 $Y=0.93
+ $X2=0.717 $Y2=0.575
r85 19 42 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.02 $X2=0.69
+ $Y2=1.935
r86 19 21 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=0.69 $Y=2.02
+ $X2=0.69 $Y2=2.815
r87 18 42 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.85 $X2=0.69
+ $Y2=1.935
r88 17 18 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=0.69 $Y=1.65 $X2=0.69
+ $Y2=1.85
r89 16 40 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.565
+ $X2=0.24 $Y2=1.48
r90 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.69 $Y2=1.65
r91 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.355 $Y2=1.565
r92 14 39 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=0.355 $Y=1.055
+ $X2=0.24 $Y2=1.18
r93 13 44 4.36636 $w=2.5e-07 $l=1.02e-07 $layer=LI1_cond $X=0.615 $Y=1.055
+ $X2=0.717 $Y2=1.055
r94 13 14 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=1.055
+ $X2=0.355 $Y2=1.055
r95 4 46 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.015
r96 4 33 400 $w=1.7e-07 $l=1.06737e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.835
r97 3 42 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r98 3 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r99 2 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.595
+ $Y=0.45 $X2=1.735 $Y2=0.595
r100 1 44 182 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.45 $X2=0.715 $Y2=1.065
r101 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.45 $X2=0.715 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%A_509_392# 1 2 3 4 5 6 21 23 24 27 29 33 37
+ 39 41 42 45 47 49 51 53 55 61 64
c103 41 0 1.12995e-19 $X=6.93 $Y=2.12
r104 57 59 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=4.76 $Y=2.375
+ $X2=4.76 $Y2=2.435
r105 55 57 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=4.76 $Y=2.085
+ $X2=4.76 $Y2=2.375
r106 49 66 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=2.12 $X2=7.88
+ $Y2=2.035
r107 49 51 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.88 $Y=2.12
+ $X2=7.88 $Y2=2.815
r108 48 63 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=2.035
+ $X2=6.93 $Y2=2.035
r109 47 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.715 $Y=2.035
+ $X2=7.88 $Y2=2.035
r110 47 48 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.715 $Y=2.035
+ $X2=7.095 $Y2=2.035
r111 43 64 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.955 $Y=2.46
+ $X2=6.93 $Y2=2.375
r112 43 45 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=6.955 $Y=2.46
+ $X2=6.955 $Y2=2.465
r113 42 64 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=2.29
+ $X2=6.93 $Y2=2.375
r114 41 63 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=2.12 $X2=6.93
+ $Y2=2.035
r115 41 42 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=6.93 $Y=2.12
+ $X2=6.93 $Y2=2.29
r116 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=2.375
+ $X2=5.95 $Y2=2.375
r117 39 64 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=2.375
+ $X2=6.93 $Y2=2.375
r118 39 40 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.765 $Y=2.375
+ $X2=6.115 $Y2=2.375
r119 35 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=2.46
+ $X2=5.95 $Y2=2.375
r120 35 37 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.95 $Y=2.46
+ $X2=5.95 $Y2=2.815
r121 34 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=2.375
+ $X2=4.76 $Y2=2.375
r122 33 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=2.375
+ $X2=5.95 $Y2=2.375
r123 33 34 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.785 $Y=2.375
+ $X2=4.925 $Y2=2.375
r124 31 59 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=4.76 $Y=2.46
+ $X2=4.76 $Y2=2.435
r125 31 32 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.76 $Y=2.46
+ $X2=4.76 $Y2=2.905
r126 30 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.99
+ $X2=3.69 $Y2=2.99
r127 29 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.595 $Y=2.99
+ $X2=4.76 $Y2=2.905
r128 29 30 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.595 $Y=2.99
+ $X2=3.855 $Y2=2.99
r129 25 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.905
+ $X2=3.69 $Y2=2.99
r130 25 27 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.69 $Y=2.905
+ $X2=3.69 $Y2=2.405
r131 23 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=2.99
+ $X2=3.69 $Y2=2.99
r132 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.525 $Y=2.99
+ $X2=2.855 $Y2=2.99
r133 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.69 $Y=2.905
+ $X2=2.855 $Y2=2.99
r134 19 21 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.69 $Y=2.905
+ $X2=2.69 $Y2=2.405
r135 6 66 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.96 $X2=7.88 $Y2=2.115
r136 6 51 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.96 $X2=7.88 $Y2=2.815
r137 5 63 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=6.78
+ $Y=1.96 $X2=6.93 $Y2=2.085
r138 5 45 300 $w=1.7e-07 $l=5.7513e-07 $layer=licon1_PDIFF $count=2 $X=6.78
+ $Y=1.96 $X2=6.93 $Y2=2.465
r139 4 61 600 $w=1.7e-07 $l=4.84226e-07 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.96 $X2=5.95 $Y2=2.375
r140 4 37 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.96 $X2=5.95 $Y2=2.815
r141 3 59 300 $w=1.7e-07 $l=5.94874e-07 $layer=licon1_PDIFF $count=2 $X=4.49
+ $Y=1.96 $X2=4.76 $Y2=2.435
r142 3 55 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.49
+ $Y=1.96 $X2=4.76 $Y2=2.085
r143 2 27 300 $w=1.7e-07 $l=5.35747e-07 $layer=licon1_PDIFF $count=2 $X=3.49
+ $Y=1.96 $X2=3.69 $Y2=2.405
r144 1 21 300 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_PDIFF $count=2 $X=2.545
+ $Y=1.96 $X2=2.69 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%VGND 1 2 3 4 5 16 18 22 26 29 32 40 41 42 44
+ 49 61 70 71 77 80 83
c89 71 0 6.39601e-20 $X=7.92 $Y=0
c90 40 0 1.36109e-20 $X=4.585 $Y=0
c91 32 0 1.9667e-19 $X=7.365 $Y=0.755
c92 1 0 3.13945e-19 $X=0.135 $Y=0.45
r93 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r94 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r95 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r96 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 71 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r98 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r99 68 83 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=7.545 $Y=0 $X2=7.367
+ $Y2=0
r100 68 70 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=0
+ $X2=7.92 $Y2=0
r101 67 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r102 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r103 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r104 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r105 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r106 61 83 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.19 $Y=0 $X2=7.367
+ $Y2=0
r107 61 66 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.19 $Y=0 $X2=6.96
+ $Y2=0
r108 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r109 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r110 57 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r111 56 59 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r112 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r113 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.235
+ $Y2=0
r114 54 56 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r115 53 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r116 53 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r117 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r118 50 77 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.195
+ $Y2=0
r119 50 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.68
+ $Y2=0
r120 49 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.235
+ $Y2=0
r121 49 52 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.68
+ $Y2=0
r122 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r123 48 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r124 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r125 45 74 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r126 45 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r127 44 77 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.195
+ $Y2=0
r128 44 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r129 42 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r130 42 57 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r131 40 59 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.56
+ $Y2=0
r132 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.67
+ $Y2=0
r133 39 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=5.04 $Y2=0
r134 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.67
+ $Y2=0
r135 30 83 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.367 $Y=0.085
+ $X2=7.367 $Y2=0
r136 30 32 21.7503 $w=3.53e-07 $l=6.7e-07 $layer=LI1_cond $X=7.367 $Y=0.085
+ $X2=7.367 $Y2=0.755
r137 29 35 9.29238 $w=1.83e-07 $l=1.55e-07 $layer=LI1_cond $X=4.67 $Y=0.847
+ $X2=4.515 $Y2=0.847
r138 28 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0
r139 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0.755
r140 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0
r141 24 26 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0.675
r142 20 77 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0
r143 20 22 14.3353 $w=4.08e-07 $l=5.1e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.595
r144 16 74 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r145 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.595
r146 5 32 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=7.215
+ $Y=0.61 $X2=7.365 $Y2=0.755
r147 4 35 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.695 $X2=4.515 $Y2=0.845
r148 3 26 91 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=2 $X=2.025
+ $Y=0.45 $X2=2.235 $Y2=0.675
r149 2 22 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.45 $X2=1.195 $Y2=0.595
r150 1 18 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.45 $X2=0.28 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%A_587_110# 1 2 9 12
c23 9 0 1.22971e-19 $X=4.015 $Y=0.84
r24 12 14 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.075 $Y=0.705
+ $X2=3.075 $Y2=0.84
r25 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0.84
+ $X2=3.075 $Y2=0.84
r26 7 9 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.24 $Y=0.84
+ $X2=4.015 $Y2=0.84
r27 2 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.695 $X2=4.015 $Y2=0.84
r28 1 12 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=2.935
+ $Y=0.55 $X2=3.075 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%A_992_122# 1 2 3 12 14 15 19 20 21 24
r48 22 24 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=7.88 $Y=1.1
+ $X2=7.88 $Y2=0.755
r49 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.715 $Y=1.185
+ $X2=7.88 $Y2=1.1
r50 20 21 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.715 $Y=1.185
+ $X2=6.99 $Y2=1.185
r51 17 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.865 $Y=1.1
+ $X2=6.99 $Y2=1.185
r52 17 19 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=6.865 $Y=1.1
+ $X2=6.865 $Y2=0.755
r53 16 19 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=6.865 $Y=0.425
+ $X2=6.865 $Y2=0.755
r54 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.74 $Y=0.34
+ $X2=6.865 $Y2=0.425
r55 14 15 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=6.74 $Y=0.34
+ $X2=5.19 $Y2=0.34
r56 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.065 $Y=0.425
+ $X2=5.19 $Y2=0.34
r57 10 12 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.065 $Y=0.425
+ $X2=5.065 $Y2=0.765
r58 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.61 $X2=7.88 $Y2=0.755
r59 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.61 $X2=6.905 $Y2=0.755
r60 1 12 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=4.96
+ $Y=0.61 $X2=5.105 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_4%A_1079_122# 1 2 7 13 16
c21 16 0 1.65419e-19 $X=6.395 $Y=0.76
c22 13 0 2.77406e-20 $X=5.535 $Y=0.765
c23 7 0 1.13206e-20 $X=6.31 $Y=0.68
r24 8 13 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.62 $Y=0.68
+ $X2=5.495 $Y2=0.68
r25 7 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.31 $Y=0.68
+ $X2=6.435 $Y2=0.68
r26 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.31 $Y=0.68 $X2=5.62
+ $Y2=0.68
r27 2 16 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=6.255
+ $Y=0.61 $X2=6.395 $Y2=0.76
r28 1 13 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.61 $X2=5.535 $Y2=0.765
.ends

