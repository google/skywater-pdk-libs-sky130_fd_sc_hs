# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__dlrbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.260000 0.835000 1.900000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.565000 0.350000 7.115000 1.050000 ;
        RECT 6.690000 1.720000 7.115000 2.850000 ;
        RECT 6.945000 1.050000 7.115000 1.720000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.195000 1.820000 8.530000 2.980000 ;
        RECT 8.245000 0.350000 8.530000 1.130000 ;
        RECT 8.360000 1.130000 8.530000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875000 1.180000 6.180000 1.550000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.260000 1.335000 1.900000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.640000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 8.830000 3.520000 ;
        RECT  1.535000 1.560000 7.080000 1.660000 ;
        RECT  5.025000 1.530000 7.080000 1.560000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.095000  0.540000 0.450000 1.090000 ;
      RECT 0.095000  1.090000 0.265000 2.070000 ;
      RECT 0.095000  2.070000 1.235000 2.240000 ;
      RECT 0.095000  2.240000 0.365000 2.980000 ;
      RECT 0.565000  2.410000 0.895000 3.245000 ;
      RECT 0.630000  0.085000 0.960000 1.090000 ;
      RECT 1.065000  2.240000 1.235000 2.730000 ;
      RECT 1.065000  2.730000 2.015000 2.900000 ;
      RECT 1.130000  0.350000 1.675000 1.090000 ;
      RECT 1.405000  2.100000 1.675000 2.220000 ;
      RECT 1.405000  2.220000 2.555000 2.390000 ;
      RECT 1.405000  2.390000 1.675000 2.560000 ;
      RECT 1.505000  1.090000 1.675000 2.100000 ;
      RECT 1.845000  0.350000 2.175000 0.780000 ;
      RECT 1.845000  0.780000 4.205000 0.950000 ;
      RECT 1.845000  0.950000 2.175000 0.960000 ;
      RECT 1.845000  0.960000 2.015000 1.720000 ;
      RECT 1.845000  1.720000 2.215000 2.050000 ;
      RECT 1.845000  2.560000 2.910000 2.730000 ;
      RECT 2.185000  1.130000 3.610000 1.300000 ;
      RECT 2.185000  1.300000 2.555000 1.550000 ;
      RECT 2.345000  0.085000 2.915000 0.600000 ;
      RECT 2.385000  1.550000 2.555000 2.220000 ;
      RECT 2.505000  2.900000 2.835000 3.245000 ;
      RECT 2.740000  1.470000 3.070000 1.800000 ;
      RECT 2.740000  1.800000 2.910000 2.560000 ;
      RECT 3.120000  1.970000 3.450000 2.140000 ;
      RECT 3.120000  2.140000 3.290000 2.905000 ;
      RECT 3.120000  2.905000 4.290000 3.075000 ;
      RECT 3.280000  1.120000 3.610000 1.130000 ;
      RECT 3.280000  1.300000 3.610000 1.450000 ;
      RECT 3.280000  1.450000 3.450000 1.970000 ;
      RECT 3.405000  0.360000 4.545000 0.610000 ;
      RECT 3.460000  2.405000 3.790000 2.735000 ;
      RECT 3.620000  1.620000 4.725000 1.790000 ;
      RECT 3.620000  1.790000 3.790000 2.405000 ;
      RECT 3.875000  0.950000 4.205000 1.450000 ;
      RECT 3.960000  2.050000 4.290000 2.905000 ;
      RECT 4.375000  0.610000 4.545000 1.220000 ;
      RECT 4.375000  1.220000 5.120000 1.550000 ;
      RECT 4.375000  1.550000 4.725000 1.620000 ;
      RECT 4.530000  1.960000 5.945000 2.290000 ;
      RECT 4.680000  2.520000 5.445000 3.245000 ;
      RECT 4.730000  0.085000 4.980000 1.030000 ;
      RECT 5.210000  0.350000 5.460000 1.050000 ;
      RECT 5.290000  1.050000 5.460000 1.720000 ;
      RECT 5.290000  1.720000 6.520000 1.890000 ;
      RECT 5.290000  1.890000 5.945000 1.960000 ;
      RECT 5.615000  2.290000 5.945000 2.850000 ;
      RECT 6.030000  0.085000 6.360000 1.010000 ;
      RECT 6.115000  2.060000 6.445000 3.245000 ;
      RECT 6.350000  1.220000 6.775000 1.550000 ;
      RECT 6.350000  1.550000 6.520000 1.720000 ;
      RECT 7.285000  0.540000 7.560000 1.300000 ;
      RECT 7.285000  1.300000 8.190000 1.630000 ;
      RECT 7.285000  1.630000 7.535000 2.780000 ;
      RECT 7.745000  0.085000 8.075000 1.130000 ;
      RECT 7.745000  1.820000 8.010000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrbn_1
END LIBRARY
