* File: sky130_fd_sc_hs__o21bai_2.spice
* Created: Tue Sep  1 20:15:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o21bai_2.pex.spice"
.subckt sky130_fd_sc_hs__o21bai_2  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_B1_N_M1012_g N_A_27_74#_M1012_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_225_74#_M1008_d N_A_27_74#_M1008_g N_Y_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1013 N_A_225_74#_M1013_d N_A_27_74#_M1013_g N_Y_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1002 N_A_225_74#_M1013_d N_A1_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1406 PD=1.09 PS=1.12 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1004 N_A_225_74#_M1004_d N_A2_M1004_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1406 PD=1.02 PS=1.12 NRD=0 NRS=4.86 M=1 R=4.93333 SA=75001.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1009 N_A_225_74#_M1004_d N_A2_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_A_225_74#_M1007_d N_A1_M1007_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_B1_N_M1003_g N_A_27_74#_M1003_s VPB PSHORT L=0.15 W=1
+ AD=0.317358 AS=0.305 PD=1.64151 PS=2.61 NRD=50.5502 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1010 N_Y_M1010_d N_A_27_74#_M1010_g N_VPWR_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.355442 PD=1.42 PS=1.83849 NRD=1.7533 NRS=14.9326 M=1 R=7.46667
+ SA=75000.9 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1010_d N_A_27_74#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2184 PD=1.42 PS=1.51 NRD=1.7533 NRS=5.2599 M=1 R=7.46667
+ SA=75001.4 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1011_s N_A1_M1000_g N_A_507_368#_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2184 AS=0.168 PD=1.51 PS=1.42 NRD=14.0658 NRS=1.7533 M=1 R=7.46667
+ SA=75001.9 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1005_d N_A2_M1005_g N_A_507_368#_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1005_d N_A2_M1006_g N_A_507_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1708 PD=1.42 PS=1.425 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_507_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.1708 PD=2.83 PS=1.425 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75003.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__o21bai_2.pxi.spice"
*
.ends
*
*
