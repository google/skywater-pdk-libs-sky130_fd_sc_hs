* File: sky130_fd_sc_hs__a32o_2.pxi.spice
* Created: Thu Aug 27 20:30:03 2020
* 
x_PM_SKY130_FD_SC_HS__A32O_2%A_45_264# N_A_45_264#_M1013_d N_A_45_264#_M1006_d
+ N_A_45_264#_c_78_n N_A_45_264#_M1010_g N_A_45_264#_M1003_g N_A_45_264#_c_79_n
+ N_A_45_264#_M1011_g N_A_45_264#_M1012_g N_A_45_264#_c_71_n N_A_45_264#_c_84_p
+ N_A_45_264#_c_114_p N_A_45_264#_c_72_n N_A_45_264#_c_86_p N_A_45_264#_c_73_n
+ N_A_45_264#_c_74_n N_A_45_264#_c_88_p N_A_45_264#_c_75_n N_A_45_264#_c_76_n
+ N_A_45_264#_c_119_p N_A_45_264#_c_110_p N_A_45_264#_c_77_n
+ PM_SKY130_FD_SC_HS__A32O_2%A_45_264#
x_PM_SKY130_FD_SC_HS__A32O_2%A3 N_A3_c_179_n N_A3_M1000_g N_A3_M1008_g A3
+ N_A3_c_181_n PM_SKY130_FD_SC_HS__A32O_2%A3
x_PM_SKY130_FD_SC_HS__A32O_2%A2 N_A2_M1007_g N_A2_c_211_n N_A2_M1002_g A2
+ N_A2_c_212_n PM_SKY130_FD_SC_HS__A32O_2%A2
x_PM_SKY130_FD_SC_HS__A32O_2%A1 N_A1_M1013_g N_A1_c_239_n N_A1_M1005_g A1
+ N_A1_c_240_n PM_SKY130_FD_SC_HS__A32O_2%A1
x_PM_SKY130_FD_SC_HS__A32O_2%B1 N_B1_M1001_g N_B1_c_270_n N_B1_M1006_g B1
+ PM_SKY130_FD_SC_HS__A32O_2%B1
x_PM_SKY130_FD_SC_HS__A32O_2%B2 N_B2_M1009_g N_B2_c_301_n N_B2_M1004_g B2
+ N_B2_c_302_n PM_SKY130_FD_SC_HS__A32O_2%B2
x_PM_SKY130_FD_SC_HS__A32O_2%VPWR N_VPWR_M1010_d N_VPWR_M1011_d N_VPWR_M1002_d
+ N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n VPWR
+ N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_321_n N_VPWR_c_330_n
+ N_VPWR_c_331_n PM_SKY130_FD_SC_HS__A32O_2%VPWR
x_PM_SKY130_FD_SC_HS__A32O_2%X N_X_M1003_s N_X_M1010_s N_X_c_376_n N_X_c_377_n X
+ N_X_c_378_n PM_SKY130_FD_SC_HS__A32O_2%X
x_PM_SKY130_FD_SC_HS__A32O_2%A_346_368# N_A_346_368#_M1000_d
+ N_A_346_368#_M1005_d N_A_346_368#_M1004_d N_A_346_368#_c_412_n
+ N_A_346_368#_c_413_n N_A_346_368#_c_421_n N_A_346_368#_c_406_n
+ N_A_346_368#_c_407_n N_A_346_368#_c_408_n N_A_346_368#_c_409_n
+ PM_SKY130_FD_SC_HS__A32O_2%A_346_368#
x_PM_SKY130_FD_SC_HS__A32O_2%VGND N_VGND_M1003_d N_VGND_M1012_d N_VGND_M1009_d
+ N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n
+ N_VGND_c_454_n VGND N_VGND_c_455_n N_VGND_c_456_n N_VGND_c_457_n
+ PM_SKY130_FD_SC_HS__A32O_2%VGND
cc_1 VNB N_A_45_264#_M1003_g 0.0282752f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_2 VNB N_A_45_264#_M1012_g 0.0244304f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.74
cc_3 VNB N_A_45_264#_c_71_n 3.74074e-19 $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.32
cc_4 VNB N_A_45_264#_c_72_n 0.00921004f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.95
cc_5 VNB N_A_45_264#_c_73_n 0.0335619f $X=-0.19 $Y=-0.245 $X2=2.775 $Y2=1.095
cc_6 VNB N_A_45_264#_c_74_n 8.19761e-19 $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.095
cc_7 VNB N_A_45_264#_c_75_n 0.00342903f $X=-0.19 $Y=-0.245 $X2=2.94 $Y2=0.515
cc_8 VNB N_A_45_264#_c_76_n 0.00395055f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.485
cc_9 VNB N_A_45_264#_c_77_n 0.0813695f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.542
cc_10 VNB N_A3_c_179_n 0.028647f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=0.37
cc_11 VNB N_A3_M1008_g 0.0265047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A3_c_181_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_13 VNB N_A2_M1007_g 0.0254275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_211_n 0.0270252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_212_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_16 VNB N_A1_M1013_g 0.0278022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_239_n 0.0250768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_240_n 0.00414591f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_19 VNB N_B1_M1001_g 0.0285948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_270_n 0.027378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB B1 0.0133269f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_22 VNB N_B2_M1009_g 0.0298505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B2_c_301_n 0.0612826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B2_c_302_n 0.00521402f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_25 VNB N_VPWR_c_321_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_376_n 0.00240426f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_27 VNB N_X_c_377_n 0.00136575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_378_n 0.00120578f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.74
cc_29 VNB N_VGND_c_449_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.32
cc_30 VNB N_VGND_c_450_n 0.0482617f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_31 VNB N_VGND_c_451_n 0.0209012f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_32 VNB N_VGND_c_452_n 0.0099193f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.74
cc_33 VNB N_VGND_c_453_n 0.0128247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_454_n 0.040801f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.32
cc_35 VNB N_VGND_c_455_n 0.0715204f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.95
cc_36 VNB N_VGND_c_456_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_457_n 0.292107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_45_264#_c_78_n 0.0170313f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_39 VPB N_A_45_264#_c_79_n 0.0165063f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_40 VPB N_A_45_264#_c_71_n 0.00759736f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.32
cc_41 VPB N_A_45_264#_c_72_n 0.00345923f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=1.95
cc_42 VPB N_A_45_264#_c_77_n 0.0138672f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.542
cc_43 VPB N_A3_c_179_n 0.0277757f $X=-0.19 $Y=1.66 $X2=2.735 $Y2=0.37
cc_44 VPB N_A3_c_181_n 0.00305163f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_45 VPB N_A2_c_211_n 0.0282648f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A2_c_212_n 0.00245998f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_47 VPB N_A1_c_239_n 0.0270253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A1_c_240_n 0.00372419f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_49 VPB N_B1_c_270_n 0.0254564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB B1 0.00583682f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_51 VPB N_B2_c_301_n 0.0272365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_B2_c_302_n 0.00778791f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_53 VPB N_VPWR_c_322_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.32
cc_54 VPB N_VPWR_c_323_n 0.0216926f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_55 VPB N_VPWR_c_324_n 0.0145913f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_56 VPB N_VPWR_c_325_n 0.0176638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_326_n 0.0206218f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=2.405
cc_58 VPB N_VPWR_c_327_n 0.0219379f $X=-0.19 $Y=1.66 $X2=2.775 $Y2=1.095
cc_59 VPB N_VPWR_c_328_n 0.0429452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_321_n 0.0818269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_330_n 0.00786036f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.65
cc_62 VPB N_VPWR_c_331_n 0.00728331f $X=-0.19 $Y=1.66 $X2=3.54 $Y2=2.065
cc_63 VPB X 0.00134143f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_64 VPB N_X_c_378_n 8.17493e-19 $X=-0.19 $Y=1.66 $X2=1 $Y2=0.74
cc_65 VPB N_A_346_368#_c_406_n 0.0206603f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_66 VPB N_A_346_368#_c_407_n 0.00350307f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.32
cc_67 VPB N_A_346_368#_c_408_n 0.0366229f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_346_368#_c_409_n 0.00312598f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=2.405
cc_69 N_A_45_264#_c_79_n N_A3_c_179_n 0.0177676f $X=0.955 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_70 N_A_45_264#_c_84_p N_A3_c_179_n 0.00173009f $X=1.105 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_45_264#_c_72_n N_A3_c_179_n 0.00609036f $X=1.19 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_45_264#_c_86_p N_A3_c_179_n 0.00358106f $X=1.19 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_73 N_A_45_264#_c_73_n N_A3_c_179_n 0.0012572f $X=2.775 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_74 N_A_45_264#_c_88_p N_A3_c_179_n 0.0161704f $X=3.375 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_75 N_A_45_264#_c_77_n N_A3_c_179_n 0.00991742f $X=0.955 $Y=1.542 $X2=-0.19
+ $Y2=-0.245
cc_76 N_A_45_264#_M1012_g N_A3_M1008_g 0.016139f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_45_264#_c_72_n N_A3_M1008_g 0.00314558f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_78 N_A_45_264#_c_73_n N_A3_M1008_g 0.0157478f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_79 N_A_45_264#_c_72_n N_A3_c_181_n 0.0327294f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_80 N_A_45_264#_c_73_n N_A3_c_181_n 0.0247243f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_81 N_A_45_264#_c_88_p N_A3_c_181_n 0.0215605f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_82 N_A_45_264#_c_73_n N_A2_M1007_g 0.0154058f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_45_264#_c_73_n N_A2_c_211_n 0.00126003f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_84 N_A_45_264#_c_88_p N_A2_c_211_n 0.0124205f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_45_264#_c_73_n N_A2_c_212_n 0.0247243f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_86 N_A_45_264#_c_88_p N_A2_c_212_n 0.0226548f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_87 N_A_45_264#_c_73_n N_A1_M1013_g 0.0161075f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_88 N_A_45_264#_c_75_n N_A1_M1013_g 0.00449149f $X=2.94 $Y=0.515 $X2=0 $Y2=0
cc_89 N_A_45_264#_c_73_n N_A1_c_239_n 0.00136523f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_90 N_A_45_264#_c_88_p N_A1_c_239_n 0.0123616f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_91 N_A_45_264#_c_73_n N_A1_c_240_n 0.030842f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_92 N_A_45_264#_c_88_p N_A1_c_240_n 0.0270914f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_45_264#_c_73_n N_B1_M1001_g 0.00292704f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_94 N_A_45_264#_c_75_n N_B1_M1001_g 0.0044057f $X=2.94 $Y=0.515 $X2=0 $Y2=0
cc_95 N_A_45_264#_c_88_p N_B1_c_270_n 0.0150046f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_45_264#_c_110_p N_B1_c_270_n 6.22879e-19 $X=3.54 $Y=2.065 $X2=0 $Y2=0
cc_97 N_A_45_264#_c_88_p B1 0.0139779f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_45_264#_c_110_p B1 0.0271963f $X=3.54 $Y=2.065 $X2=0 $Y2=0
cc_99 N_A_45_264#_c_71_n N_VPWR_M1010_d 0.0209621f $X=0.31 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_45_264#_c_114_p N_VPWR_M1010_d 0.00950867f $X=0.395 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_101 N_A_45_264#_c_84_p N_VPWR_M1011_d 0.00572185f $X=1.105 $Y=2.405 $X2=0
+ $Y2=0
cc_102 N_A_45_264#_c_72_n N_VPWR_M1011_d 0.00325404f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_103 N_A_45_264#_c_86_p N_VPWR_M1011_d 0.0054773f $X=1.19 $Y=2.32 $X2=0 $Y2=0
cc_104 N_A_45_264#_c_88_p N_VPWR_M1011_d 0.0132222f $X=3.375 $Y=2.035 $X2=0
+ $Y2=0
cc_105 N_A_45_264#_c_119_p N_VPWR_M1011_d 0.00295949f $X=1.19 $Y=2.035 $X2=0
+ $Y2=0
cc_106 N_A_45_264#_c_88_p N_VPWR_M1002_d 0.0159615f $X=3.375 $Y=2.035 $X2=0
+ $Y2=0
cc_107 N_A_45_264#_c_78_n N_VPWR_c_323_n 0.0111655f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_A_45_264#_c_79_n N_VPWR_c_323_n 0.00131191f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_45_264#_c_84_p N_VPWR_c_323_n 0.00100103f $X=1.105 $Y=2.405 $X2=0
+ $Y2=0
cc_110 N_A_45_264#_c_114_p N_VPWR_c_323_n 0.0129795f $X=0.395 $Y=2.405 $X2=0
+ $Y2=0
cc_111 N_A_45_264#_c_79_n N_VPWR_c_324_n 0.00889766f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_A_45_264#_c_84_p N_VPWR_c_324_n 0.0148723f $X=1.105 $Y=2.405 $X2=0
+ $Y2=0
cc_113 N_A_45_264#_c_88_p N_VPWR_c_324_n 0.00802589f $X=3.375 $Y=2.035 $X2=0
+ $Y2=0
cc_114 N_A_45_264#_c_78_n N_VPWR_c_326_n 0.00413917f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_45_264#_c_79_n N_VPWR_c_326_n 0.00461464f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A_45_264#_c_78_n N_VPWR_c_321_n 0.00414505f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_45_264#_c_79_n N_VPWR_c_321_n 0.00469135f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_45_264#_c_84_p N_VPWR_c_321_n 0.0214206f $X=1.105 $Y=2.405 $X2=0
+ $Y2=0
cc_119 N_A_45_264#_c_114_p N_VPWR_c_321_n 6.15054e-19 $X=0.395 $Y=2.405 $X2=0
+ $Y2=0
cc_120 N_A_45_264#_c_84_p N_X_M1010_s 0.00557733f $X=1.105 $Y=2.405 $X2=0 $Y2=0
cc_121 N_A_45_264#_M1003_g N_X_c_376_n 0.00868565f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A_45_264#_M1012_g N_X_c_376_n 0.0107619f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_45_264#_M1003_g N_X_c_377_n 0.00327408f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_45_264#_M1012_g N_X_c_377_n 0.00221233f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_45_264#_c_74_n N_X_c_377_n 0.00969158f $X=1.275 $Y=1.095 $X2=0 $Y2=0
cc_126 N_A_45_264#_c_78_n X 0.00438198f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_45_264#_c_79_n X 0.0051073f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A_45_264#_c_71_n X 0.013316f $X=0.31 $Y=2.32 $X2=0 $Y2=0
cc_129 N_A_45_264#_c_84_p X 0.0197697f $X=1.105 $Y=2.405 $X2=0 $Y2=0
cc_130 N_A_45_264#_c_86_p X 0.00219866f $X=1.19 $Y=2.32 $X2=0 $Y2=0
cc_131 N_A_45_264#_c_119_p X 0.0141517f $X=1.19 $Y=2.035 $X2=0 $Y2=0
cc_132 N_A_45_264#_c_77_n X 0.00523067f $X=0.955 $Y=1.542 $X2=0 $Y2=0
cc_133 N_A_45_264#_M1003_g N_X_c_378_n 0.00286404f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_45_264#_c_79_n N_X_c_378_n 0.00125633f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_45_264#_M1012_g N_X_c_378_n 0.00323488f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_45_264#_c_71_n N_X_c_378_n 0.00576043f $X=0.31 $Y=2.32 $X2=0 $Y2=0
cc_137 N_A_45_264#_c_72_n N_X_c_378_n 0.0564948f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_138 N_A_45_264#_c_76_n N_X_c_378_n 0.0239356f $X=0.39 $Y=1.485 $X2=0 $Y2=0
cc_139 N_A_45_264#_c_77_n N_X_c_378_n 0.0232034f $X=0.955 $Y=1.542 $X2=0 $Y2=0
cc_140 N_A_45_264#_c_88_p N_A_346_368#_M1000_d 0.00907415f $X=3.375 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_141 N_A_45_264#_c_88_p N_A_346_368#_M1005_d 0.00907415f $X=3.375 $Y=2.035
+ $X2=0 $Y2=0
cc_142 N_A_45_264#_c_88_p N_A_346_368#_c_412_n 0.0506274f $X=3.375 $Y=2.035
+ $X2=0 $Y2=0
cc_143 N_A_45_264#_c_88_p N_A_346_368#_c_413_n 0.0173337f $X=3.375 $Y=2.035
+ $X2=0 $Y2=0
cc_144 N_A_45_264#_c_110_p N_A_346_368#_c_406_n 0.0237369f $X=3.54 $Y=2.065
+ $X2=0 $Y2=0
cc_145 N_A_45_264#_c_79_n N_A_346_368#_c_409_n 7.6973e-19 $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_146 N_A_45_264#_c_84_p N_A_346_368#_c_409_n 0.00701023f $X=1.105 $Y=2.405
+ $X2=0 $Y2=0
cc_147 N_A_45_264#_c_86_p N_A_346_368#_c_409_n 0.00110648f $X=1.19 $Y=2.32 $X2=0
+ $Y2=0
cc_148 N_A_45_264#_c_88_p N_A_346_368#_c_409_n 0.017089f $X=3.375 $Y=2.035 $X2=0
+ $Y2=0
cc_149 N_A_45_264#_c_73_n N_VGND_M1012_d 0.00551645f $X=2.775 $Y=1.095 $X2=0
+ $Y2=0
cc_150 N_A_45_264#_c_74_n N_VGND_M1012_d 0.00421237f $X=1.275 $Y=1.095 $X2=0
+ $Y2=0
cc_151 N_A_45_264#_M1003_g N_VGND_c_450_n 0.019585f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_45_264#_c_76_n N_VGND_c_450_n 0.0176651f $X=0.39 $Y=1.485 $X2=0 $Y2=0
cc_153 N_A_45_264#_c_77_n N_VGND_c_450_n 0.00169922f $X=0.955 $Y=1.542 $X2=0
+ $Y2=0
cc_154 N_A_45_264#_M1003_g N_VGND_c_451_n 0.00439591f $X=0.56 $Y=0.74 $X2=0
+ $Y2=0
cc_155 N_A_45_264#_M1012_g N_VGND_c_451_n 0.00451103f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_45_264#_M1012_g N_VGND_c_452_n 0.00798291f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_45_264#_c_73_n N_VGND_c_452_n 0.0194082f $X=2.775 $Y=1.095 $X2=0
+ $Y2=0
cc_158 N_A_45_264#_c_74_n N_VGND_c_452_n 0.0080244f $X=1.275 $Y=1.095 $X2=0
+ $Y2=0
cc_159 N_A_45_264#_c_75_n N_VGND_c_455_n 0.0146357f $X=2.94 $Y=0.515 $X2=0 $Y2=0
cc_160 N_A_45_264#_M1003_g N_VGND_c_457_n 0.00842009f $X=0.56 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_45_264#_M1012_g N_VGND_c_457_n 0.00878376f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_45_264#_c_75_n N_VGND_c_457_n 0.0121141f $X=2.94 $Y=0.515 $X2=0 $Y2=0
cc_163 N_A_45_264#_c_73_n A_355_74# 0.0048076f $X=2.775 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_45_264#_c_73_n A_433_74# 0.0120044f $X=2.775 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A3_M1008_g N_A2_M1007_g 0.0395125f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A3_c_179_n N_A2_c_211_n 0.0669304f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A3_c_181_n N_A2_c_211_n 0.00178024f $X=1.61 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A3_c_179_n N_A2_c_212_n 0.00137132f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A3_c_181_n N_A2_c_212_n 0.0249837f $X=1.61 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A3_c_179_n N_VPWR_c_324_n 0.00561023f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A3_c_179_n N_VPWR_c_327_n 0.00481995f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A3_c_179_n N_VPWR_c_321_n 0.00508379f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A3_M1008_g N_X_c_376_n 8.11115e-19 $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A3_c_179_n N_A_346_368#_c_409_n 0.00956742f $X=1.655 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A3_M1008_g N_VGND_c_452_n 0.0168903f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A3_M1008_g N_VGND_c_455_n 0.00461464f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A3_M1008_g N_VGND_c_457_n 0.00911119f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A2_M1007_g N_A1_M1013_g 0.0343511f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A2_c_211_n N_A1_c_239_n 0.0407341f $X=2.105 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A2_c_212_n N_A1_c_239_n 6.37986e-19 $X=2.18 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A2_c_211_n N_A1_c_240_n 0.00233311f $X=2.105 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A2_c_212_n N_A1_c_240_n 0.0334556f $X=2.18 $Y=1.515 $X2=0 $Y2=0
cc_183 N_A2_c_211_n N_VPWR_c_325_n 0.00583349f $X=2.105 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A2_c_211_n N_VPWR_c_327_n 0.00481995f $X=2.105 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A2_c_211_n N_VPWR_c_321_n 0.00508379f $X=2.105 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A2_c_211_n N_A_346_368#_c_412_n 0.0126982f $X=2.105 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A2_c_211_n N_A_346_368#_c_421_n 7.55911e-19 $X=2.105 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A2_c_211_n N_A_346_368#_c_409_n 0.00703033f $X=2.105 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A2_M1007_g N_VGND_c_455_n 0.00461464f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A2_M1007_g N_VGND_c_457_n 0.0091028f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A1_M1013_g N_B1_M1001_g 0.0261158f $X=2.66 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_c_239_n N_B1_c_270_n 0.0452967f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A1_c_240_n N_B1_c_270_n 7.86772e-19 $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A1_c_239_n B1 0.00161275f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A1_c_240_n B1 0.0266982f $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A1_c_239_n N_VPWR_c_325_n 0.00373226f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A1_c_239_n N_VPWR_c_328_n 0.00451897f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A1_c_239_n N_VPWR_c_321_n 0.00457541f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A1_c_239_n N_A_346_368#_c_412_n 0.0126982f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A1_c_239_n N_A_346_368#_c_413_n 4.27055e-19 $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A1_c_239_n N_A_346_368#_c_421_n 0.00754046f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A1_c_239_n N_A_346_368#_c_407_n 0.00178875f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A1_c_239_n N_A_346_368#_c_409_n 7.45827e-19 $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A1_M1013_g N_VGND_c_455_n 0.00461464f $X=2.66 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A1_M1013_g N_VGND_c_457_n 0.00911823f $X=2.66 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B1_M1001_g N_B2_M1009_g 0.0306717f $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B1_c_270_n N_B2_c_301_n 0.0493737f $X=3.265 $Y=1.765 $X2=0 $Y2=0
cc_208 B1 N_B2_c_301_n 0.00400625f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_209 N_B1_M1001_g N_B2_c_302_n 2.13129e-19 $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B1_c_270_n N_B2_c_302_n 2.84591e-19 $X=3.265 $Y=1.765 $X2=0 $Y2=0
cc_211 B1 N_B2_c_302_n 0.0354768f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_212 N_B1_c_270_n N_VPWR_c_328_n 7.44201e-19 $X=3.265 $Y=1.765 $X2=0 $Y2=0
cc_213 N_B1_c_270_n N_A_346_368#_c_413_n 0.00184286f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_B1_c_270_n N_A_346_368#_c_421_n 0.00672358f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_B1_c_270_n N_A_346_368#_c_406_n 0.00990262f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_216 N_B1_c_270_n N_A_346_368#_c_407_n 0.00114023f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_217 N_B1_c_270_n N_A_346_368#_c_408_n 7.60962e-19 $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_B1_M1001_g N_VGND_c_454_n 0.00407036f $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_219 N_B1_M1001_g N_VGND_c_455_n 0.00461464f $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_220 N_B1_M1001_g N_VGND_c_457_n 0.00911823f $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B2_c_301_n N_VPWR_c_328_n 7.44201e-19 $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_222 N_B2_c_301_n N_A_346_368#_c_421_n 5.78806e-19 $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_B2_c_301_n N_A_346_368#_c_406_n 0.0115629f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_224 N_B2_c_301_n N_A_346_368#_c_408_n 0.01907f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_225 N_B2_c_302_n N_A_346_368#_c_408_n 0.0258667f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_226 N_B2_M1009_g N_VGND_c_454_n 0.0240799f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B2_c_301_n N_VGND_c_454_n 0.00285025f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_228 N_B2_c_302_n N_VGND_c_454_n 0.0254821f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_229 N_B2_M1009_g N_VGND_c_455_n 0.00383152f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B2_M1009_g N_VGND_c_457_n 0.00758792f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_231 N_VPWR_M1002_d N_A_346_368#_c_412_n 0.0130432f $X=2.18 $Y=1.84 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_325_n N_A_346_368#_c_412_n 0.0307535f $X=2.46 $Y=2.715 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_325_n N_A_346_368#_c_421_n 0.0171894f $X=2.46 $Y=2.715 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_328_n N_A_346_368#_c_406_n 0.0667586f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_321_n N_A_346_368#_c_406_n 0.0380121f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_325_n N_A_346_368#_c_407_n 0.0119784f $X=2.46 $Y=2.715 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_328_n N_A_346_368#_c_407_n 0.0236566f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_321_n N_A_346_368#_c_407_n 0.0128296f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_324_n N_A_346_368#_c_409_n 0.0137045f $X=1.305 $Y=2.825 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_325_n N_A_346_368#_c_409_n 0.0148394f $X=2.46 $Y=2.715 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_327_n N_A_346_368#_c_409_n 0.0096394f $X=2.265 $Y=3.33 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_321_n N_A_346_368#_c_409_n 0.011097f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_243 N_X_c_376_n N_VGND_c_450_n 0.0322525f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_244 N_X_c_376_n N_VGND_c_451_n 0.0153382f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_245 N_X_c_376_n N_VGND_c_452_n 0.0294488f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_246 N_X_c_376_n N_VGND_c_457_n 0.0117503f $X=0.78 $Y=0.495 $X2=0 $Y2=0
