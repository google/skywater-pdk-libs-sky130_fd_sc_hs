* File: sky130_fd_sc_hs__sdfxtp_1.spice
* Created: Tue Sep  1 20:23:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfxtp_1.pex.spice"
.subckt sky130_fd_sc_hs__sdfxtp_1  VNB VPB SCE D SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_SCE_M1006_g N_A_35_74#_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.07455 AS=0.1197 PD=0.775 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1014 A_223_74# N_A_35_74#_M1014_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.07455 PD=0.66 PS=0.775 NRD=18.564 NRS=21.42 M=1 R=2.8
+ SA=75000.7 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_301_74#_M1015_d N_D_M1015_g A_223_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.12495 AS=0.0504 PD=1.015 PS=0.66 NRD=48.564 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1026 A_450_74# N_SCE_M1026_g N_A_301_74#_M1015_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.12495 PD=0.66 PS=1.015 NRD=18.564 NRS=41.424 M=1 R=2.8
+ SA=75001.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_SCD_M1024_g A_450_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0504 PD=0.796552 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_630_74#_M1003_d N_CLK_M1003_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.154634 PD=2.05 PS=1.40345 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_A_828_74#_M1013_d N_A_630_74#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.2109 PD=2.01 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_1018_100#_M1007_d N_A_630_74#_M1007_g N_A_301_74#_M1007_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=0.95 PS=1.37 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1028 A_1154_100# N_A_828_74#_M1028_g N_A_1018_100#_M1007_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08925 AS=0.1113 PD=0.845 PS=0.95 NRD=45 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75004.1 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_1239_74#_M1018_g A_1154_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.174387 AS=0.08925 PD=1.19505 PS=0.845 NRD=102.912 NRS=45 M=1 R=2.8
+ SA=75001.4 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1010 N_A_1239_74#_M1010_d N_A_1018_100#_M1010_g N_VGND_M1018_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.078375 AS=0.228363 PD=0.835 PS=1.56495 NRD=1.08 NRS=72 M=1
+ R=3.66667 SA=75001.9 SB=75002.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_1520_74#_M1000_d N_A_828_74#_M1000_g N_A_1239_74#_M1010_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.182747 AS=0.078375 PD=1.40619 PS=0.835 NRD=89.448 NRS=0 M=1
+ R=3.66667 SA=75002.3 SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1017 A_1688_100# N_A_630_74#_M1017_g N_A_1520_74#_M1000_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.139553 PD=0.66 PS=1.07381 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75003.5 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_1736_74#_M1004_g A_1688_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.140462 AS=0.0504 PD=1.07814 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.9
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 N_A_1736_74#_M1008_d N_A_1520_74#_M1008_g N_VGND_M1004_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.183938 PD=1.63 PS=1.41186 NRD=0 NRS=15.264 M=1
+ R=3.66667 SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1012 N_Q_M1012_d N_A_1736_74#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.1998 PD=2.03 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_VPWR_M1019_d N_SCE_M1019_g N_A_35_74#_M1019_s VPB PSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1888 PD=0.99 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1020 A_238_464# N_SCE_M1020_g N_VPWR_M1019_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1005 N_A_301_74#_M1005_d N_D_M1005_g A_238_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1009 A_412_464# N_A_35_74#_M1009_g N_A_301_74#_M1005_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1248 AS=0.096 PD=1.03 PS=0.94 NRD=43.0839 NRS=3.0732 M=1 R=4.26667
+ SA=75001.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1022 N_VPWR_M1022_d N_SCD_M1022_g A_412_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.176582 AS=0.1248 PD=1.22182 PS=1.03 NRD=55.3964 NRS=43.0839 M=1 R=4.26667
+ SA=75002.1 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1025 N_A_630_74#_M1025_d N_CLK_M1025_g N_VPWR_M1022_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.309018 PD=2.83 PS=2.13818 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75001.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1027 N_A_828_74#_M1027_d N_A_630_74#_M1027_g N_VPWR_M1027_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.532 PD=2.83 PS=3.19 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75000.4 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1031 N_A_1018_100#_M1031_d N_A_828_74#_M1031_g N_A_301_74#_M1031_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1239 PD=0.77 PS=1.43 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1029 A_1202_508# N_A_630_74#_M1029_g N_A_1018_100#_M1031_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0525 AS=0.0735 PD=0.67 PS=0.77 NRD=32.8202 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_1239_74#_M1002_g A_1202_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.1232 AS=0.0525 PD=1.01333 PS=0.67 NRD=46.886 NRS=32.8202 M=1 R=2.8
+ SA=75001.1 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1023 N_A_1239_74#_M1023_d N_A_1018_100#_M1023_g N_VPWR_M1002_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2331 AS=0.2464 PD=1.395 PS=2.02667 NRD=0 NRS=55.8889 M=1
+ R=5.6 SA=75001 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1030 N_A_1520_74#_M1030_d N_A_630_74#_M1030_g N_A_1239_74#_M1023_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2618 AS=0.2331 PD=1.86 PS=1.395 NRD=22.261 NRS=58.6272 M=1
+ R=5.6 SA=75001.7 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1016 A_1688_508# N_A_828_74#_M1016_g N_A_1520_74#_M1030_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1309 PD=0.69 PS=0.93 NRD=37.5088 NRS=84.4145 M=1 R=2.8
+ SA=75003.1 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_1736_74#_M1001_g A_1688_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.1204 AS=0.0567 PD=0.956667 PS=0.69 NRD=60.9715 NRS=37.5088 M=1 R=2.8
+ SA=75003.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1021 N_A_1736_74#_M1021_d N_A_1520_74#_M1021_g N_VPWR_M1001_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2478 AS=0.2408 PD=2.27 PS=1.91333 NRD=2.3443 NRS=43.3794
+ M=1 R=5.6 SA=75002.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_Q_M1011_d N_A_1736_74#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3248 AS=0.3304 PD=2.82 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=21.2412 P=26.56
c_122 VNB 0 2.44411e-19 $X=0 $Y=0
c_223 VPB 0 3.2853e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__sdfxtp_1.pxi.spice"
*
.ends
*
*
