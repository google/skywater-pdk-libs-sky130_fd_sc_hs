* NGSPICE file created from sky130_fd_sc_hs__o41a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR B1 a_428_368# VPB pshort w=1e+06u l=150000u
+  ad=1.7526e+12p pd=1.002e+07u as=4.554e+11p ps=3.08e+06u
M1001 a_200_368# A2 a_116_368# VPB pshort w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=3.024e+11p ps=2.78e+06u
M1002 X a_428_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1003 VPWR a_428_368# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=6.364e+11p pd=6.16e+06u as=1.2691e+12p ps=9.35e+06u
M1005 X a_428_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_116_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_428_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_428_368# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1010 a_428_368# A4 a_314_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1011 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_314_368# A3 a_200_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

