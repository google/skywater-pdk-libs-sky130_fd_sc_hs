* File: sky130_fd_sc_hs__o221a_1.pxi.spice
* Created: Tue Sep  1 20:15:26 2020
* 
x_PM_SKY130_FD_SC_HS__O221A_1%A_83_264# N_A_83_264#_M1005_d N_A_83_264#_M1006_d
+ N_A_83_264#_M1011_d N_A_83_264#_c_73_n N_A_83_264#_M1009_g N_A_83_264#_M1003_g
+ N_A_83_264#_c_79_n N_A_83_264#_c_80_n N_A_83_264#_c_134_p N_A_83_264#_c_81_n
+ N_A_83_264#_c_103_p N_A_83_264#_c_82_n N_A_83_264#_c_75_n N_A_83_264#_c_76_n
+ N_A_83_264#_c_84_n N_A_83_264#_c_77_n N_A_83_264#_c_85_n
+ PM_SKY130_FD_SC_HS__O221A_1%A_83_264#
x_PM_SKY130_FD_SC_HS__O221A_1%A1 N_A1_M1002_g N_A1_c_163_n N_A1_M1004_g A1
+ PM_SKY130_FD_SC_HS__O221A_1%A1
x_PM_SKY130_FD_SC_HS__O221A_1%A2 N_A2_M1000_g N_A2_c_196_n N_A2_M1006_g A2
+ PM_SKY130_FD_SC_HS__O221A_1%A2
x_PM_SKY130_FD_SC_HS__O221A_1%B2 N_B2_c_227_n N_B2_c_228_n N_B2_M1010_g
+ N_B2_c_229_n N_B2_c_230_n N_B2_c_231_n N_B2_M1001_g B2
+ PM_SKY130_FD_SC_HS__O221A_1%B2
x_PM_SKY130_FD_SC_HS__O221A_1%B1 N_B1_c_272_n N_B1_M1008_g N_B1_M1007_g B1
+ N_B1_c_271_n PM_SKY130_FD_SC_HS__O221A_1%B1
x_PM_SKY130_FD_SC_HS__O221A_1%C1 N_C1_c_305_n N_C1_M1005_g N_C1_c_310_n
+ N_C1_M1011_g C1 C1 N_C1_c_307_n N_C1_c_308_n PM_SKY130_FD_SC_HS__O221A_1%C1
x_PM_SKY130_FD_SC_HS__O221A_1%X N_X_M1003_s N_X_M1009_s N_X_c_345_n N_X_c_346_n
+ N_X_c_342_n X X N_X_c_344_n X PM_SKY130_FD_SC_HS__O221A_1%X
x_PM_SKY130_FD_SC_HS__O221A_1%VPWR N_VPWR_M1009_d N_VPWR_M1008_d N_VPWR_c_366_n
+ N_VPWR_c_367_n VPWR N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_365_n
+ N_VPWR_c_371_n N_VPWR_c_372_n PM_SKY130_FD_SC_HS__O221A_1%VPWR
x_PM_SKY130_FD_SC_HS__O221A_1%VGND N_VGND_M1003_d N_VGND_M1000_d N_VGND_c_408_n
+ N_VGND_c_409_n N_VGND_c_410_n N_VGND_c_411_n VGND N_VGND_c_412_n
+ N_VGND_c_413_n N_VGND_c_414_n PM_SKY130_FD_SC_HS__O221A_1%VGND
x_PM_SKY130_FD_SC_HS__O221A_1%A_245_94# N_A_245_94#_M1002_d N_A_245_94#_M1001_d
+ N_A_245_94#_c_452_n N_A_245_94#_c_453_n N_A_245_94#_c_454_n
+ N_A_245_94#_c_471_n PM_SKY130_FD_SC_HS__O221A_1%A_245_94#
x_PM_SKY130_FD_SC_HS__O221A_1%A_456_74# N_A_456_74#_M1001_s N_A_456_74#_M1007_d
+ N_A_456_74#_c_488_n N_A_456_74#_c_489_n N_A_456_74#_c_490_n
+ N_A_456_74#_c_498_n PM_SKY130_FD_SC_HS__O221A_1%A_456_74#
cc_1 VNB N_A_83_264#_c_73_n 0.0390543f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_83_264#_M1003_g 0.0301825f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.74
cc_3 VNB N_A_83_264#_c_75_n 0.0333404f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=1.96
cc_4 VNB N_A_83_264#_c_76_n 0.00390048f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.485
cc_5 VNB N_A_83_264#_c_77_n 0.0271336f $X=-0.19 $Y=-0.245 $X2=3.935 $Y2=0.525
cc_6 VNB N_A1_M1002_g 0.0313341f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=1.96
cc_7 VNB N_A1_c_163_n 0.0198093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A1 0.00325184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_M1000_g 0.0316315f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=1.96
cc_10 VNB N_A2_c_196_n 0.0165935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A2 0.00299813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B2_c_227_n 0.0282098f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.96
cc_13 VNB N_B2_c_228_n 0.00280391f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=1.96
cc_14 VNB N_B2_c_229_n 0.0194238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_c_230_n 0.0199768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B2_c_231_n 0.0194669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB B2 0.00444804f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB N_B1_M1007_g 0.0359828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB B1 0.00248798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_271_n 0.026171f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_21 VNB N_C1_c_305_n 0.0265844f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.96
cc_22 VNB C1 0.00795525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_c_307_n 0.0237545f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.74
cc_24 VNB N_C1_c_308_n 0.0218548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_342_n 0.0250068f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.74
cc_26 VNB X 0.0145164f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.65
cc_27 VNB N_X_c_344_n 0.0273847f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=2.815
cc_28 VNB N_VPWR_c_365_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_408_n 0.0236354f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_30 VNB N_VGND_c_409_n 0.016373f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.65
cc_31 VNB N_VGND_c_410_n 0.01947f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.035
cc_32 VNB N_VGND_c_411_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=2.13
cc_33 VNB N_VGND_c_412_n 0.0587016f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=1.96
cc_34 VNB N_VGND_c_413_n 0.267882f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.485
cc_35 VNB N_VGND_c_414_n 0.0272997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_245_94#_c_452_n 0.00327588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_245_94#_c_453_n 0.0216121f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_38 VNB N_A_245_94#_c_454_n 0.00406832f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_39 VNB N_A_456_74#_c_488_n 0.00465728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_456_74#_c_489_n 0.00490525f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_41 VNB N_A_456_74#_c_490_n 0.00489174f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_42 VPB N_A_83_264#_c_73_n 0.0303537f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_43 VPB N_A_83_264#_c_79_n 0.00289739f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_44 VPB N_A_83_264#_c_80_n 0.0106319f $X=-0.19 $Y=1.66 $X2=1.725 $Y2=2.035
cc_45 VPB N_A_83_264#_c_81_n 0.00299332f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=2.815
cc_46 VPB N_A_83_264#_c_82_n 0.0350163f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.815
cc_47 VPB N_A_83_264#_c_75_n 0.0141695f $X=-0.19 $Y=1.66 $X2=4.12 $Y2=1.96
cc_48 VPB N_A_83_264#_c_84_n 0.0037217f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=2.115
cc_49 VPB N_A_83_264#_c_85_n 0.0106334f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.125
cc_50 VPB N_A1_c_163_n 0.0386029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB A1 0.00138199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A2_c_196_n 0.0343567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB A2 0.00174709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_B2_c_228_n 0.0365408f $X=-0.19 $Y=1.66 $X2=3.89 $Y2=1.96
cc_55 VPB B2 0.00311741f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_56 VPB N_B1_c_272_n 0.0202109f $X=-0.19 $Y=1.66 $X2=3.725 $Y2=0.37
cc_57 VPB B1 0.00304223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B1_c_271_n 0.0307107f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_59 VPB N_C1_c_305_n 0.0261123f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.96
cc_60 VPB N_C1_c_310_n 0.0230811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB C1 0.00314059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_X_c_345_n 0.0118064f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_63 VPB N_X_c_346_n 0.0405221f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.32
cc_64 VPB N_X_c_342_n 0.00737672f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=0.74
cc_65 VPB N_VPWR_c_366_n 0.0105397f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_66 VPB N_VPWR_c_367_n 0.0119956f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=0.74
cc_67 VPB N_VPWR_c_368_n 0.0546548f $X=-0.19 $Y=1.66 $X2=1.725 $Y2=2.035
cc_68 VPB N_VPWR_c_369_n 0.0191515f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.815
cc_69 VPB N_VPWR_c_365_n 0.0948595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_371_n 0.0285033f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.485
cc_71 VPB N_VPWR_c_372_n 0.015951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 N_A_83_264#_c_73_n N_A1_M1002_g 0.00601582f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_83_264#_M1003_g N_A1_M1002_g 0.0202137f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_83_264#_c_76_n N_A1_M1002_g 8.05667e-19 $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_75 N_A_83_264#_c_73_n N_A1_c_163_n 0.0319309f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_83_264#_c_79_n N_A1_c_163_n 0.00408813f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_77 N_A_83_264#_c_80_n N_A1_c_163_n 0.0179803f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_78 N_A_83_264#_c_81_n N_A1_c_163_n 0.00285895f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_79 N_A_83_264#_c_76_n N_A1_c_163_n 7.10742e-19 $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_80 N_A_83_264#_c_73_n A1 7.26157e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_83_264#_c_80_n A1 0.0242115f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_82 N_A_83_264#_c_76_n A1 0.0202352f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_83 N_A_83_264#_c_80_n N_A2_c_196_n 0.012228f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_84 N_A_83_264#_c_81_n N_A2_c_196_n 0.0160851f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_85 N_A_83_264#_c_84_n N_A2_c_196_n 0.00466649f $X=1.89 $Y=2.115 $X2=0 $Y2=0
cc_86 N_A_83_264#_c_80_n A2 0.0115269f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_87 N_A_83_264#_c_84_n A2 0.0151122f $X=1.89 $Y=2.115 $X2=0 $Y2=0
cc_88 N_A_83_264#_c_81_n N_B2_c_228_n 0.0229846f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_89 N_A_83_264#_c_103_p N_B2_c_228_n 0.0202163f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_90 N_A_83_264#_c_84_n N_B2_c_228_n 3.13634e-19 $X=1.89 $Y=2.115 $X2=0 $Y2=0
cc_91 N_A_83_264#_c_103_p B2 0.0391746f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_92 N_A_83_264#_c_103_p N_B1_c_272_n 0.0206639f $X=3.875 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_83_264#_c_103_p B1 0.0239398f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_94 N_A_83_264#_c_103_p N_B1_c_271_n 0.0022741f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_95 N_A_83_264#_c_103_p N_C1_c_305_n 0.00150877f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_96 N_A_83_264#_c_103_p N_C1_c_310_n 0.0154515f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_97 N_A_83_264#_c_82_n N_C1_c_310_n 0.0144886f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_98 N_A_83_264#_c_75_n N_C1_c_310_n 8.62041e-19 $X=4.12 $Y=1.96 $X2=0 $Y2=0
cc_99 N_A_83_264#_c_85_n N_C1_c_310_n 9.50925e-19 $X=4.04 $Y=2.125 $X2=0 $Y2=0
cc_100 N_A_83_264#_c_103_p C1 0.0242925f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_101 N_A_83_264#_c_75_n C1 0.0429988f $X=4.12 $Y=1.96 $X2=0 $Y2=0
cc_102 N_A_83_264#_c_77_n C1 0.00409207f $X=3.935 $Y=0.525 $X2=0 $Y2=0
cc_103 N_A_83_264#_c_75_n N_C1_c_307_n 0.020227f $X=4.12 $Y=1.96 $X2=0 $Y2=0
cc_104 N_A_83_264#_c_77_n N_C1_c_307_n 0.00420768f $X=3.935 $Y=0.525 $X2=0 $Y2=0
cc_105 N_A_83_264#_c_75_n N_C1_c_308_n 0.00352354f $X=4.12 $Y=1.96 $X2=0 $Y2=0
cc_106 N_A_83_264#_c_77_n N_C1_c_308_n 0.0114582f $X=3.935 $Y=0.525 $X2=0 $Y2=0
cc_107 N_A_83_264#_c_73_n N_X_c_345_n 0.00349474f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_83_264#_c_79_n N_X_c_345_n 0.00559275f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_109 N_A_83_264#_c_73_n N_X_c_346_n 0.0181528f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_83_264#_c_73_n N_X_c_342_n 0.010641f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_83_264#_M1003_g N_X_c_342_n 0.00457487f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_83_264#_c_79_n N_X_c_342_n 0.00566753f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_113 N_A_83_264#_c_76_n N_X_c_342_n 0.0248004f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_114 N_A_83_264#_c_73_n X 0.00220539f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_83_264#_M1003_g X 0.00285885f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_83_264#_c_76_n X 0.00479823f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_117 N_A_83_264#_M1003_g N_X_c_344_n 0.00787957f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_83_264#_c_79_n N_VPWR_M1009_d 0.00239213f $X=0.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_83_264#_c_80_n N_VPWR_M1009_d 0.00902889f $X=1.725 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_83_264#_c_134_p N_VPWR_M1009_d 0.0045173f $X=0.785 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_83_264#_c_103_p N_VPWR_M1008_d 0.0254954f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_122 N_A_83_264#_c_73_n N_VPWR_c_366_n 0.0113032f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_83_264#_c_80_n N_VPWR_c_366_n 0.0222558f $X=1.725 $Y=2.035 $X2=0
+ $Y2=0
cc_124 N_A_83_264#_c_134_p N_VPWR_c_366_n 0.00933174f $X=0.785 $Y=2.035 $X2=0
+ $Y2=0
cc_125 N_A_83_264#_c_81_n N_VPWR_c_366_n 0.0183153f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_126 N_A_83_264#_c_103_p N_VPWR_c_367_n 0.0617178f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_127 N_A_83_264#_c_82_n N_VPWR_c_367_n 0.0263973f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_128 N_A_83_264#_c_81_n N_VPWR_c_368_n 0.0145938f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_129 N_A_83_264#_c_82_n N_VPWR_c_369_n 0.0145938f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_130 N_A_83_264#_c_73_n N_VPWR_c_365_n 0.00863959f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_83_264#_c_81_n N_VPWR_c_365_n 0.0120466f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_132 N_A_83_264#_c_82_n N_VPWR_c_365_n 0.0120466f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_133 N_A_83_264#_c_73_n N_VPWR_c_371_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A_83_264#_c_80_n A_264_392# 0.00595227f $X=1.725 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A_83_264#_c_103_p A_462_392# 0.0153213f $X=3.875 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_83_264#_c_73_n N_VGND_c_408_n 7.25643e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_83_264#_M1003_g N_VGND_c_408_n 0.00946427f $X=0.57 $Y=0.74 $X2=0
+ $Y2=0
cc_138 N_A_83_264#_c_76_n N_VGND_c_408_n 0.00762027f $X=0.62 $Y=1.485 $X2=0
+ $Y2=0
cc_139 N_A_83_264#_c_77_n N_VGND_c_412_n 0.018459f $X=3.935 $Y=0.525 $X2=0 $Y2=0
cc_140 N_A_83_264#_M1003_g N_VGND_c_413_n 0.00828947f $X=0.57 $Y=0.74 $X2=0
+ $Y2=0
cc_141 N_A_83_264#_c_77_n N_VGND_c_413_n 0.0158482f $X=3.935 $Y=0.525 $X2=0
+ $Y2=0
cc_142 N_A_83_264#_M1003_g N_VGND_c_414_n 0.00434272f $X=0.57 $Y=0.74 $X2=0
+ $Y2=0
cc_143 N_A_83_264#_c_80_n N_A_245_94#_c_453_n 9.96677e-19 $X=1.725 $Y=2.035
+ $X2=0 $Y2=0
cc_144 N_A_83_264#_c_84_n N_A_245_94#_c_453_n 0.00484566f $X=1.89 $Y=2.115 $X2=0
+ $Y2=0
cc_145 N_A_83_264#_M1003_g N_A_245_94#_c_454_n 6.79941e-19 $X=0.57 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_83_264#_c_80_n N_A_245_94#_c_454_n 0.00633136f $X=1.725 $Y=2.035
+ $X2=0 $Y2=0
cc_147 N_A_83_264#_c_77_n N_A_456_74#_c_489_n 0.00313012f $X=3.935 $Y=0.525
+ $X2=0 $Y2=0
cc_148 N_A1_M1002_g N_A2_M1000_g 0.0248377f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_149 N_A1_c_163_n N_A2_c_196_n 0.078759f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_150 A1 N_A2_c_196_n 4.11485e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A1_c_163_n A2 0.00200717f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_152 A1 A2 0.020843f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A1_c_163_n N_VPWR_c_366_n 0.0145947f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_154 N_A1_c_163_n N_VPWR_c_368_n 0.00461464f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_155 N_A1_c_163_n N_VPWR_c_365_n 0.00911633f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_156 N_A1_M1002_g N_VGND_c_408_n 0.00744236f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_157 A1 N_VGND_c_408_n 6.86881e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A1_M1002_g N_VGND_c_409_n 6.44645e-19 $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_159 N_A1_M1002_g N_VGND_c_410_n 0.00485498f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_160 N_A1_M1002_g N_VGND_c_413_n 0.00514438f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_161 N_A1_M1002_g N_A_245_94#_c_452_n 0.00748716f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_162 N_A1_M1002_g N_A_245_94#_c_454_n 0.0062738f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_163 N_A1_c_163_n N_A_245_94#_c_454_n 8.5326e-19 $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_164 A1 N_A_245_94#_c_454_n 0.0112432f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A2_c_196_n N_B2_c_227_n 0.0181454f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_166 A2 N_B2_c_227_n 4.19338e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A2_c_196_n N_B2_c_228_n 0.0210241f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_168 N_A2_M1000_g N_B2_c_230_n 0.011086f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_169 N_A2_c_196_n B2 4.16298e-19 $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_170 A2 B2 0.0197629f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A2_c_196_n N_VPWR_c_368_n 0.00445602f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_172 N_A2_c_196_n N_VPWR_c_365_n 0.00859212f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_173 N_A2_M1000_g N_VGND_c_409_n 0.0122599f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_174 N_A2_M1000_g N_VGND_c_410_n 0.00421418f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_175 N_A2_M1000_g N_VGND_c_413_n 0.00432128f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_176 N_A2_M1000_g N_A_245_94#_c_452_n 0.00350341f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_177 N_A2_M1000_g N_A_245_94#_c_453_n 0.0153207f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_178 N_A2_c_196_n N_A_245_94#_c_453_n 0.00411453f $X=1.665 $Y=1.885 $X2=0
+ $Y2=0
cc_179 A2 N_A_245_94#_c_453_n 0.0250329f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A2_M1000_g N_A_456_74#_c_488_n 0.00116577f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_181 N_A2_M1000_g N_A_456_74#_c_490_n 3.62451e-19 $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_182 N_B2_c_228_n N_B1_c_272_n 0.0332151f $X=2.235 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_183 N_B2_c_227_n N_B1_M1007_g 0.00510377f $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_184 N_B2_c_231_n N_B1_M1007_g 0.0275047f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_185 B2 N_B1_M1007_g 2.17586e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_186 N_B2_c_227_n B1 2.35705e-19 $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_187 B2 B1 0.0260436f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_188 N_B2_c_227_n N_B1_c_271_n 0.00387701f $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_189 N_B2_c_228_n N_B1_c_271_n 0.0117842f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_190 N_B2_c_229_n N_B1_c_271_n 0.00238913f $X=2.645 $Y=1.175 $X2=0 $Y2=0
cc_191 B2 N_B1_c_271_n 0.00649914f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_192 N_B2_c_228_n N_VPWR_c_367_n 0.00352484f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_193 N_B2_c_228_n N_VPWR_c_368_n 0.00461464f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_194 N_B2_c_228_n N_VPWR_c_365_n 0.00911823f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_195 N_B2_c_231_n N_VGND_c_409_n 7.83914e-19 $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_196 N_B2_c_231_n N_VGND_c_412_n 0.00278271f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_197 N_B2_c_231_n N_VGND_c_413_n 0.00358525f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_198 N_B2_c_227_n N_A_245_94#_c_453_n 0.0063832f $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_199 N_B2_c_229_n N_A_245_94#_c_453_n 0.0178297f $X=2.645 $Y=1.175 $X2=0 $Y2=0
cc_200 N_B2_c_230_n N_A_245_94#_c_453_n 0.0118983f $X=2.475 $Y=1.175 $X2=0 $Y2=0
cc_201 B2 N_A_245_94#_c_453_n 0.0457618f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_202 N_B2_c_229_n N_A_245_94#_c_471_n 5.20128e-19 $X=2.645 $Y=1.175 $X2=0
+ $Y2=0
cc_203 N_B2_c_231_n N_A_245_94#_c_471_n 0.0123389f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_204 N_B2_c_230_n N_A_456_74#_c_488_n 0.00812328f $X=2.475 $Y=1.175 $X2=0
+ $Y2=0
cc_205 N_B2_c_231_n N_A_456_74#_c_489_n 0.0133401f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_206 B1 N_C1_c_305_n 4.13026e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_207 N_B1_c_271_n N_C1_c_305_n 0.0178735f $X=3.09 $Y=1.625 $X2=0 $Y2=0
cc_208 N_B1_M1007_g C1 0.00496568f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_209 B1 C1 0.0208926f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_210 N_B1_c_271_n C1 0.00207338f $X=3.09 $Y=1.625 $X2=0 $Y2=0
cc_211 N_B1_M1007_g N_C1_c_307_n 0.0147786f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_212 N_B1_M1007_g N_C1_c_308_n 0.017212f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_213 N_B1_c_272_n N_VPWR_c_367_n 0.0213519f $X=2.805 $Y=1.885 $X2=0 $Y2=0
cc_214 N_B1_c_272_n N_VPWR_c_368_n 0.00413917f $X=2.805 $Y=1.885 $X2=0 $Y2=0
cc_215 N_B1_c_272_n N_VPWR_c_365_n 0.00818781f $X=2.805 $Y=1.885 $X2=0 $Y2=0
cc_216 N_B1_M1007_g N_VGND_c_412_n 0.00278271f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_217 N_B1_M1007_g N_VGND_c_413_n 0.00354237f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_218 N_B1_M1007_g N_A_245_94#_c_453_n 0.00516704f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_219 B1 N_A_245_94#_c_453_n 0.0140154f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_220 N_B1_c_271_n N_A_245_94#_c_453_n 0.00698857f $X=3.09 $Y=1.625 $X2=0 $Y2=0
cc_221 N_B1_M1007_g N_A_245_94#_c_471_n 0.0084974f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_222 N_B1_M1007_g N_A_456_74#_c_489_n 0.0133206f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_223 N_C1_c_310_n N_VPWR_c_367_n 0.0185782f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_224 N_C1_c_310_n N_VPWR_c_369_n 0.00445602f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_225 N_C1_c_310_n N_VPWR_c_365_n 0.00865213f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_226 N_C1_c_308_n N_VGND_c_412_n 0.00430908f $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_227 N_C1_c_308_n N_VGND_c_413_n 0.00821503f $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_228 C1 N_A_245_94#_c_453_n 0.00728498f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_229 N_C1_c_308_n N_A_245_94#_c_471_n 6.13134e-19 $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_230 N_C1_c_308_n N_A_456_74#_c_489_n 0.00735461f $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_231 C1 N_A_456_74#_c_498_n 0.00723658f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_232 N_C1_c_307_n N_A_456_74#_c_498_n 4.53017e-19 $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_233 N_C1_c_308_n N_A_456_74#_c_498_n 0.0059147f $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_234 N_X_c_346_n N_VPWR_c_366_n 0.0422702f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_235 N_X_c_346_n N_VPWR_c_365_n 0.0120466f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_236 N_X_c_346_n N_VPWR_c_371_n 0.0145938f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_237 N_X_c_344_n N_VGND_c_408_n 0.0317414f $X=0.355 $Y=0.515 $X2=0 $Y2=0
cc_238 N_X_c_344_n N_VGND_c_413_n 0.0147684f $X=0.355 $Y=0.515 $X2=0 $Y2=0
cc_239 N_X_c_344_n N_VGND_c_414_n 0.0179105f $X=0.355 $Y=0.515 $X2=0 $Y2=0
cc_240 N_VGND_c_408_n N_A_245_94#_c_452_n 0.0243787f $X=0.855 $Y=0.515 $X2=0
+ $Y2=0
cc_241 N_VGND_c_409_n N_A_245_94#_c_452_n 0.0191765f $X=1.865 $Y=0.735 $X2=0
+ $Y2=0
cc_242 N_VGND_c_410_n N_A_245_94#_c_452_n 0.0103491f $X=1.7 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_413_n N_A_245_94#_c_452_n 0.0113354f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_244 N_VGND_c_409_n N_A_245_94#_c_453_n 0.0244412f $X=1.865 $Y=0.735 $X2=0
+ $Y2=0
cc_245 N_VGND_c_408_n N_A_245_94#_c_454_n 0.00156673f $X=0.855 $Y=0.515 $X2=0
+ $Y2=0
cc_246 N_VGND_c_409_n N_A_456_74#_c_488_n 0.0346871f $X=1.865 $Y=0.735 $X2=0
+ $Y2=0
cc_247 N_VGND_c_412_n N_A_456_74#_c_489_n 0.0664804f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_413_n N_A_456_74#_c_489_n 0.0369159f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_409_n N_A_456_74#_c_490_n 0.0121618f $X=1.865 $Y=0.735 $X2=0
+ $Y2=0
cc_250 N_VGND_c_412_n N_A_456_74#_c_490_n 0.0236697f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_251 N_VGND_c_413_n N_A_456_74#_c_490_n 0.0128321f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_252 N_A_245_94#_c_453_n N_A_456_74#_c_488_n 0.0258597f $X=2.77 $Y=1.195 $X2=0
+ $Y2=0
cc_253 N_A_245_94#_M1001_d N_A_456_74#_c_489_n 0.00176461f $X=2.795 $Y=0.37
+ $X2=0 $Y2=0
cc_254 N_A_245_94#_c_471_n N_A_456_74#_c_489_n 0.016064f $X=2.935 $Y=0.81 $X2=0
+ $Y2=0
