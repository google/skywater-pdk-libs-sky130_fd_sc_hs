* File: sky130_fd_sc_hs__buf_8.pxi.spice
* Created: Thu Aug 27 20:34:42 2020
* 
x_PM_SKY130_FD_SC_HS__BUF_8%A N_A_M1001_g N_A_c_108_n N_A_M1004_g N_A_c_109_n
+ N_A_M1005_g N_A_M1015_g N_A_M1019_g N_A_c_110_n N_A_M1007_g A A A N_A_c_106_n
+ N_A_c_107_n PM_SKY130_FD_SC_HS__BUF_8%A
x_PM_SKY130_FD_SC_HS__BUF_8%A_27_74# N_A_27_74#_M1001_d N_A_27_74#_M1015_d
+ N_A_27_74#_M1004_d N_A_27_74#_M1005_d N_A_27_74#_M1000_g N_A_27_74#_c_187_n
+ N_A_27_74#_M1003_g N_A_27_74#_M1002_g N_A_27_74#_c_188_n N_A_27_74#_M1008_g
+ N_A_27_74#_M1006_g N_A_27_74#_c_189_n N_A_27_74#_M1009_g N_A_27_74#_M1012_g
+ N_A_27_74#_c_190_n N_A_27_74#_M1010_g N_A_27_74#_M1016_g N_A_27_74#_c_191_n
+ N_A_27_74#_M1011_g N_A_27_74#_M1017_g N_A_27_74#_c_192_n N_A_27_74#_M1013_g
+ N_A_27_74#_c_193_n N_A_27_74#_M1014_g N_A_27_74#_M1020_g N_A_27_74#_M1021_g
+ N_A_27_74#_c_194_n N_A_27_74#_M1018_g N_A_27_74#_c_178_n N_A_27_74#_c_195_n
+ N_A_27_74#_c_196_n N_A_27_74#_c_179_n N_A_27_74#_c_180_n N_A_27_74#_c_212_n
+ N_A_27_74#_c_197_n N_A_27_74#_c_181_n N_A_27_74#_c_182_n N_A_27_74#_c_224_n
+ N_A_27_74#_c_183_n N_A_27_74#_c_248_p N_A_27_74#_c_227_n N_A_27_74#_c_184_n
+ N_A_27_74#_c_185_n N_A_27_74#_c_186_n PM_SKY130_FD_SC_HS__BUF_8%A_27_74#
x_PM_SKY130_FD_SC_HS__BUF_8%VPWR N_VPWR_M1004_s N_VPWR_M1007_s N_VPWR_M1008_s
+ N_VPWR_M1010_s N_VPWR_M1013_s N_VPWR_M1018_s N_VPWR_c_402_n N_VPWR_c_403_n
+ N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n
+ VPWR N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n N_VPWR_c_412_n
+ N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n
+ N_VPWR_c_418_n N_VPWR_c_401_n PM_SKY130_FD_SC_HS__BUF_8%VPWR
x_PM_SKY130_FD_SC_HS__BUF_8%X N_X_M1000_d N_X_M1006_d N_X_M1016_d N_X_M1020_d
+ N_X_M1003_d N_X_M1009_d N_X_M1011_d N_X_M1014_d N_X_c_490_n N_X_c_502_n
+ N_X_c_491_n N_X_c_492_n N_X_c_503_n N_X_c_504_n N_X_c_493_n N_X_c_505_n
+ N_X_c_494_n N_X_c_506_n N_X_c_495_n N_X_c_507_n N_X_c_496_n N_X_c_508_n
+ N_X_c_497_n N_X_c_498_n N_X_c_499_n N_X_c_510_n N_X_c_500_n N_X_c_511_n
+ N_X_c_501_n X X X X PM_SKY130_FD_SC_HS__BUF_8%X
x_PM_SKY130_FD_SC_HS__BUF_8%VGND N_VGND_M1001_s N_VGND_M1019_s N_VGND_M1002_s
+ N_VGND_M1012_s N_VGND_M1017_s N_VGND_M1021_s N_VGND_c_645_n N_VGND_c_646_n
+ N_VGND_c_647_n N_VGND_c_648_n N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n
+ N_VGND_c_652_n N_VGND_c_653_n N_VGND_c_654_n N_VGND_c_655_n N_VGND_c_656_n
+ N_VGND_c_657_n VGND N_VGND_c_658_n N_VGND_c_659_n N_VGND_c_660_n
+ N_VGND_c_661_n N_VGND_c_662_n N_VGND_c_663_n PM_SKY130_FD_SC_HS__BUF_8%VGND
cc_1 VNB N_A_M1001_g 0.0325279f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_M1015_g 0.0237982f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_3 VNB N_A_M1019_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_4 VNB N_A_c_106_n 0.0166485f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_5 VNB N_A_c_107_n 0.0567134f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.557
cc_6 VNB N_A_27_74#_M1000_g 0.0197781f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.35
cc_7 VNB N_A_27_74#_M1002_g 0.0212166f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A_27_74#_M1006_g 0.0217898f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_9 VNB N_A_27_74#_M1012_g 0.0225551f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_10 VNB N_A_27_74#_M1016_g 0.0225551f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_11 VNB N_A_27_74#_M1017_g 0.0225551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_M1020_g 0.0225878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_M1021_g 0.02608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_178_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_179_n 0.00351687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_180_n 0.00998227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_181_n 0.00179731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_182_n 0.0043023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_183_n 4.30857e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_184_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_185_n 0.00335789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_186_n 0.242206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_401_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_490_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_491_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.557
cc_26 VNB N_X_c_492_n 0.00140587f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_27 VNB N_X_c_493_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_494_n 0.00311987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_495_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_496_n 0.00311987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_497_n 0.0024448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_498_n 0.00141267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_499_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_500_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_501_n 0.00181295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_645_n 0.0055945f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_37 VNB N_VGND_c_646_n 0.00256838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_647_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_39 VNB N_VGND_c_648_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.557
cc_40 VNB N_VGND_c_649_n 0.00831705f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_41 VNB N_VGND_c_650_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.557
cc_42 VNB N_VGND_c_651_n 0.0551405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_652_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_44 VNB N_VGND_c_653_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_654_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_655_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.565
cc_47 VNB N_VGND_c_656_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_657_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_658_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_659_n 0.0167636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_660_n 0.0188148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_661_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_662_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_663_n 0.322609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_A_c_108_n 0.0208611f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_56 VPB N_A_c_109_n 0.0155109f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_57 VPB N_A_c_110_n 0.0158647f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_58 VPB N_A_c_106_n 0.0138362f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_59 VPB N_A_c_107_n 0.0344451f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.557
cc_60 VPB N_A_27_74#_c_187_n 0.0155806f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_61 VPB N_A_27_74#_c_188_n 0.0160039f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_62 VPB N_A_27_74#_c_189_n 0.0156201f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_63 VPB N_A_27_74#_c_190_n 0.015621f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.557
cc_64 VPB N_A_27_74#_c_191_n 0.0156201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_27_74#_c_192_n 0.0155121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_27_74#_c_193_n 0.0157041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_74#_c_194_n 0.0175368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_27_74#_c_195_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_74#_c_196_n 0.0353617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_74#_c_197_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_74#_c_183_n 0.00287436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_74#_c_186_n 0.056321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_402_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_74 VPB N_VPWR_c_403_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_404_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_76 VPB N_VPWR_c_405_n 0.00886117f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.557
cc_77 VPB N_VPWR_c_406_n 0.00891739f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.557
cc_78 VPB N_VPWR_c_407_n 0.0120875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_408_n 0.0645735f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.565
cc_80 VPB N_VPWR_c_409_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_410_n 0.0194914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_411_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_412_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_413_n 0.0195976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_414_n 0.0234893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_415_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_416_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_417_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_418_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_401_n 0.0849977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_X_c_502_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_92 VPB N_X_c_503_n 0.00209566f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_93 VPB N_X_c_504_n 0.00232642f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.557
cc_94 VPB N_X_c_505_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_X_c_506_n 0.00209566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_X_c_507_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_X_c_508_n 0.00200554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_X_c_498_n 8.47603e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_X_c_510_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_X_c_511_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB X 0.00138058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB X 0.00290135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 N_A_M1019_g N_A_27_74#_M1000_g 0.0311454f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_c_110_n N_A_27_74#_c_187_n 0.0221126f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_M1001_g N_A_27_74#_c_178_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_c_108_n N_A_27_74#_c_195_n 4.27055e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A_c_106_n N_A_27_74#_c_195_n 0.0260502f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A_c_108_n N_A_27_74#_c_196_n 0.0104891f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A_c_109_n N_A_27_74#_c_196_n 6.45594e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_M1001_g N_A_27_74#_c_179_n 0.0139147f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_M1015_g N_A_27_74#_c_179_n 0.0140682f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_c_106_n N_A_27_74#_c_179_n 0.0554204f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_113 N_A_c_107_n N_A_27_74#_c_179_n 0.00325098f $X=1.4 $Y=1.557 $X2=0 $Y2=0
cc_114 N_A_c_106_n N_A_27_74#_c_180_n 0.0216404f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A_c_108_n N_A_27_74#_c_212_n 0.0120074f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_c_109_n N_A_27_74#_c_212_n 0.0120074f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_c_106_n N_A_27_74#_c_212_n 0.0393875f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A_c_107_n N_A_27_74#_c_212_n 0.00131177f $X=1.4 $Y=1.557 $X2=0 $Y2=0
cc_119 N_A_c_108_n N_A_27_74#_c_197_n 6.45594e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_c_109_n N_A_27_74#_c_197_n 0.0103431f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_c_110_n N_A_27_74#_c_197_n 0.0104721f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_M1015_g N_A_27_74#_c_181_n 4.04737e-19 $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_M1019_g N_A_27_74#_c_181_n 3.92313e-19 $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_M1019_g N_A_27_74#_c_182_n 0.0135996f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_c_106_n N_A_27_74#_c_182_n 0.0118433f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A_c_107_n N_A_27_74#_c_182_n 9.9484e-19 $X=1.4 $Y=1.557 $X2=0 $Y2=0
cc_127 N_A_c_110_n N_A_27_74#_c_224_n 0.0133273f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A_c_106_n N_A_27_74#_c_224_n 0.00580317f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A_c_110_n N_A_27_74#_c_183_n 0.00389155f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_c_109_n N_A_27_74#_c_227_n 4.27055e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_c_110_n N_A_27_74#_c_227_n 4.27055e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A_c_106_n N_A_27_74#_c_227_n 0.0237598f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_107_n N_A_27_74#_c_227_n 0.00144162f $X=1.4 $Y=1.557 $X2=0 $Y2=0
cc_134 N_A_c_106_n N_A_27_74#_c_184_n 0.0146029f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A_c_107_n N_A_27_74#_c_184_n 0.00232957f $X=1.4 $Y=1.557 $X2=0 $Y2=0
cc_136 N_A_M1019_g N_A_27_74#_c_185_n 0.00394038f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_c_106_n N_A_27_74#_c_185_n 0.0341212f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_c_107_n N_A_27_74#_c_185_n 0.0030667f $X=1.4 $Y=1.557 $X2=0 $Y2=0
cc_139 N_A_c_106_n N_A_27_74#_c_186_n 2.37596e-19 $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A_c_107_n N_A_27_74#_c_186_n 0.0196911f $X=1.4 $Y=1.557 $X2=0 $Y2=0
cc_141 N_A_c_108_n N_VPWR_c_402_n 0.00486623f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_c_109_n N_VPWR_c_402_n 0.00486623f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_c_110_n N_VPWR_c_403_n 0.00526215f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_c_109_n N_VPWR_c_409_n 0.00445602f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_c_110_n N_VPWR_c_409_n 0.00445602f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_c_108_n N_VPWR_c_414_n 0.00445602f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_c_108_n N_VPWR_c_401_n 0.008611f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_c_109_n N_VPWR_c_401_n 0.00857589f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_c_110_n N_VPWR_c_401_n 0.00857673f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A_M1001_g N_VGND_c_645_n 0.0136079f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_M1015_g N_VGND_c_645_n 0.00238937f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_M1015_g N_VGND_c_646_n 4.78024e-19 $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_M1019_g N_VGND_c_646_n 0.010688f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_M1001_g N_VGND_c_658_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_M1015_g N_VGND_c_659_n 0.00461464f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_M1019_g N_VGND_c_659_n 0.00383152f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_M1001_g N_VGND_c_663_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A_M1015_g N_VGND_c_663_n 0.00907982f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_M1019_g N_VGND_c_663_n 0.0075754f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_27_74#_c_212_n N_VPWR_M1004_s 0.00408911f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_27_74#_c_224_n N_VPWR_M1007_s 0.00499186f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_162 N_A_27_74#_c_183_n N_VPWR_M1007_s 0.00160462f $X=1.685 $Y=1.95 $X2=0
+ $Y2=0
cc_163 N_A_27_74#_c_196_n N_VPWR_c_402_n 0.0449718f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_164 N_A_27_74#_c_212_n N_VPWR_c_402_n 0.0136682f $X=1.02 $Y=2.035 $X2=0 $Y2=0
cc_165 N_A_27_74#_c_197_n N_VPWR_c_402_n 0.0449718f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_166 N_A_27_74#_c_187_n N_VPWR_c_403_n 0.0105202f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A_27_74#_c_188_n N_VPWR_c_403_n 7.03309e-19 $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_27_74#_c_197_n N_VPWR_c_403_n 0.0462948f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_169 N_A_27_74#_c_224_n N_VPWR_c_403_n 0.0154457f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_170 N_A_27_74#_c_248_p N_VPWR_c_403_n 5.27207e-19 $X=4.64 $Y=1.465 $X2=0
+ $Y2=0
cc_171 N_A_27_74#_c_188_n N_VPWR_c_404_n 0.00646055f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A_27_74#_c_189_n N_VPWR_c_404_n 0.00750878f $X=2.86 $Y=1.765 $X2=0
+ $Y2=0
cc_173 N_A_27_74#_c_190_n N_VPWR_c_405_n 0.00646055f $X=3.31 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A_27_74#_c_191_n N_VPWR_c_405_n 0.00750878f $X=3.81 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A_27_74#_c_192_n N_VPWR_c_406_n 0.00641457f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_A_27_74#_c_193_n N_VPWR_c_406_n 0.00381884f $X=4.745 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A_27_74#_c_194_n N_VPWR_c_408_n 0.00999852f $X=5.21 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A_27_74#_c_197_n N_VPWR_c_409_n 0.014552f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_179 N_A_27_74#_c_187_n N_VPWR_c_410_n 0.00413917f $X=1.86 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A_27_74#_c_188_n N_VPWR_c_410_n 0.00445602f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_27_74#_c_189_n N_VPWR_c_411_n 0.00445602f $X=2.86 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_27_74#_c_190_n N_VPWR_c_411_n 0.00445602f $X=3.31 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_27_74#_c_191_n N_VPWR_c_412_n 0.00445602f $X=3.81 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A_27_74#_c_192_n N_VPWR_c_412_n 0.00445602f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_27_74#_c_193_n N_VPWR_c_413_n 0.00461464f $X=4.745 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_27_74#_c_194_n N_VPWR_c_413_n 0.00439937f $X=5.21 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_27_74#_c_196_n N_VPWR_c_414_n 0.0145938f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_188 N_A_27_74#_c_187_n N_VPWR_c_401_n 0.00818187f $X=1.86 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A_27_74#_c_188_n N_VPWR_c_401_n 0.00858511f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A_27_74#_c_189_n N_VPWR_c_401_n 0.00857378f $X=2.86 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A_27_74#_c_190_n N_VPWR_c_401_n 0.0085805f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_27_74#_c_191_n N_VPWR_c_401_n 0.00857378f $X=3.81 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_27_74#_c_192_n N_VPWR_c_401_n 0.00857917f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_A_27_74#_c_193_n N_VPWR_c_401_n 0.00908413f $X=4.745 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_27_74#_c_194_n N_VPWR_c_401_n 0.00843023f $X=5.21 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_27_74#_c_196_n N_VPWR_c_401_n 0.0120466f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_197 N_A_27_74#_c_197_n N_VPWR_c_401_n 0.0119791f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_198 N_A_27_74#_M1000_g N_X_c_490_n 3.92313e-19 $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_27_74#_M1002_g N_X_c_490_n 3.92313e-19 $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_27_74#_c_187_n N_X_c_502_n 0.00543866f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_27_74#_c_188_n N_X_c_502_n 0.0127211f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_27_74#_c_189_n N_X_c_502_n 7.39949e-19 $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_27_74#_M1002_g N_X_c_491_n 0.0128315f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_27_74#_M1006_g N_X_c_491_n 0.0115433f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_27_74#_c_248_p N_X_c_491_n 0.0500092f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_206 N_A_27_74#_c_186_n N_X_c_491_n 0.00387558f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_207 N_A_27_74#_c_248_p N_X_c_492_n 0.0143381f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_208 N_A_27_74#_c_185_n N_X_c_492_n 0.00455444f $X=1.685 $Y=1.095 $X2=0 $Y2=0
cc_209 N_A_27_74#_c_186_n N_X_c_492_n 0.00232957f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_210 N_A_27_74#_c_188_n N_X_c_503_n 0.0122806f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A_27_74#_c_189_n N_X_c_503_n 0.0122806f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A_27_74#_c_248_p N_X_c_503_n 0.0455181f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_213 N_A_27_74#_c_186_n N_X_c_503_n 0.00875137f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_214 N_A_27_74#_c_187_n N_X_c_504_n 0.00108872f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A_27_74#_c_188_n N_X_c_504_n 9.20137e-19 $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A_27_74#_c_183_n N_X_c_504_n 0.00293378f $X=1.685 $Y=1.95 $X2=0 $Y2=0
cc_217 N_A_27_74#_c_248_p N_X_c_504_n 0.0277622f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_218 N_A_27_74#_c_186_n N_X_c_504_n 0.00825852f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_219 N_A_27_74#_M1002_g N_X_c_493_n 8.71574e-19 $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_27_74#_M1006_g N_X_c_493_n 0.0089455f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_27_74#_M1012_g N_X_c_493_n 0.00916694f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_27_74#_M1016_g N_X_c_493_n 6.18925e-19 $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_27_74#_c_188_n N_X_c_505_n 6.39139e-19 $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A_27_74#_c_189_n N_X_c_505_n 0.0121613f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A_27_74#_c_190_n N_X_c_505_n 0.0127555f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A_27_74#_c_191_n N_X_c_505_n 7.39949e-19 $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A_27_74#_M1012_g N_X_c_494_n 0.0118691f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_27_74#_M1016_g N_X_c_494_n 0.0118691f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A_27_74#_c_248_p N_X_c_494_n 0.0493541f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_230 N_A_27_74#_c_186_n N_X_c_494_n 0.00552382f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_231 N_A_27_74#_c_190_n N_X_c_506_n 0.0122806f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_27_74#_c_191_n N_X_c_506_n 0.0122806f $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_27_74#_c_248_p N_X_c_506_n 0.0455181f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_234 N_A_27_74#_c_186_n N_X_c_506_n 0.00855438f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_235 N_A_27_74#_M1012_g N_X_c_495_n 6.18925e-19 $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_27_74#_M1016_g N_X_c_495_n 0.00916694f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A_27_74#_M1017_g N_X_c_495_n 0.00916694f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_27_74#_M1020_g N_X_c_495_n 6.18925e-19 $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A_27_74#_c_190_n N_X_c_507_n 6.39139e-19 $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_27_74#_c_191_n N_X_c_507_n 0.0121613f $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_27_74#_c_192_n N_X_c_507_n 0.0127197f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_27_74#_c_193_n N_X_c_507_n 6.79477e-19 $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_27_74#_M1017_g N_X_c_496_n 0.0118691f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_27_74#_M1020_g N_X_c_496_n 0.0118144f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A_27_74#_c_248_p N_X_c_496_n 0.0490309f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_186_n N_X_c_496_n 0.00538093f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_247 N_A_27_74#_c_192_n N_X_c_508_n 0.0122025f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A_27_74#_c_193_n N_X_c_508_n 0.0135147f $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_27_74#_c_248_p N_X_c_508_n 0.0444246f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_250 N_A_27_74#_c_186_n N_X_c_508_n 0.00802155f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_251 N_A_27_74#_M1017_g N_X_c_497_n 6.18848e-19 $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_27_74#_M1020_g N_X_c_497_n 0.00918133f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_27_74#_M1021_g N_X_c_497_n 0.00768946f $X=5.195 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_27_74#_M1020_g N_X_c_498_n 0.00257778f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_27_74#_M1021_g N_X_c_498_n 0.00858408f $X=5.195 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_27_74#_c_194_n N_X_c_498_n 0.00194866f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_27_74#_c_248_p N_X_c_498_n 0.0249855f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_258 N_A_27_74#_c_186_n N_X_c_498_n 0.0369565f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_259 N_A_27_74#_M1006_g N_X_c_499_n 9.7541e-19 $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_27_74#_M1012_g N_X_c_499_n 9.7541e-19 $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_27_74#_c_248_p N_X_c_499_n 0.0276081f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_262 N_A_27_74#_c_186_n N_X_c_499_n 0.00239372f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_263 N_A_27_74#_c_189_n N_X_c_510_n 9.3899e-19 $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_27_74#_c_190_n N_X_c_510_n 9.3899e-19 $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A_27_74#_c_248_p N_X_c_510_n 0.0276943f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_266 N_A_27_74#_c_186_n N_X_c_510_n 0.00798099f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_267 N_A_27_74#_M1016_g N_X_c_500_n 9.7541e-19 $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_27_74#_M1017_g N_X_c_500_n 9.7541e-19 $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_27_74#_c_248_p N_X_c_500_n 0.0276081f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_270 N_A_27_74#_c_186_n N_X_c_500_n 0.00232957f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_271 N_A_27_74#_c_191_n N_X_c_511_n 9.3899e-19 $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A_27_74#_c_192_n N_X_c_511_n 9.3899e-19 $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_273 N_A_27_74#_c_248_p N_X_c_511_n 0.0276943f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_274 N_A_27_74#_c_186_n N_X_c_511_n 0.00792231f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_275 N_A_27_74#_M1020_g N_X_c_501_n 0.00130353f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_27_74#_M1021_g N_X_c_501_n 0.00205051f $X=5.195 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A_27_74#_c_186_n N_X_c_501_n 0.00150825f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_278 N_A_27_74#_c_193_n X 5.13605e-19 $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_279 N_A_27_74#_c_194_n X 0.00362003f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A_27_74#_c_186_n X 0.00519017f $X=5.195 $Y=1.532 $X2=0 $Y2=0
cc_281 N_A_27_74#_c_193_n X 4.30474e-19 $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_282 N_A_27_74#_c_194_n X 0.0120377f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_283 N_A_27_74#_c_179_n N_VGND_M1001_s 0.00224297f $X=1.1 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_284 N_A_27_74#_c_182_n N_VGND_M1019_s 9.61034e-19 $X=1.6 $Y=1.095 $X2=0 $Y2=0
cc_285 N_A_27_74#_c_185_n N_VGND_M1019_s 0.00130977f $X=1.685 $Y=1.095 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_178_n N_VGND_c_645_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_287 N_A_27_74#_c_179_n N_VGND_c_645_n 0.0189527f $X=1.1 $Y=1.095 $X2=0 $Y2=0
cc_288 N_A_27_74#_c_181_n N_VGND_c_645_n 0.00123668f $X=1.185 $Y=0.515 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_M1000_g N_VGND_c_646_n 0.01069f $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A_27_74#_M1002_g N_VGND_c_646_n 4.71636e-19 $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A_27_74#_c_181_n N_VGND_c_646_n 0.0182488f $X=1.185 $Y=0.515 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_c_182_n N_VGND_c_646_n 0.00731846f $X=1.6 $Y=1.095 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_248_p N_VGND_c_646_n 3.19484e-19 $X=4.64 $Y=1.465 $X2=0
+ $Y2=0
cc_294 N_A_27_74#_c_185_n N_VGND_c_646_n 0.00988848f $X=1.685 $Y=1.095 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_M1000_g N_VGND_c_647_n 4.56715e-19 $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A_27_74#_M1002_g N_VGND_c_647_n 0.00956829f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_27_74#_M1006_g N_VGND_c_647_n 0.00406778f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A_27_74#_M1012_g N_VGND_c_648_n 0.00454042f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_299 N_A_27_74#_M1016_g N_VGND_c_648_n 0.00454042f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_300 N_A_27_74#_M1017_g N_VGND_c_649_n 0.00454042f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_27_74#_M1020_g N_VGND_c_649_n 0.0045466f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_27_74#_M1021_g N_VGND_c_651_n 0.0184966f $X=5.195 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A_27_74#_M1000_g N_VGND_c_652_n 0.00383152f $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A_27_74#_M1002_g N_VGND_c_652_n 0.00383152f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A_27_74#_M1006_g N_VGND_c_654_n 0.00434272f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A_27_74#_M1012_g N_VGND_c_654_n 0.00434272f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_27_74#_M1016_g N_VGND_c_656_n 0.00434272f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A_27_74#_M1017_g N_VGND_c_656_n 0.00434272f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_178_n N_VGND_c_658_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_181_n N_VGND_c_659_n 0.00749631f $X=1.185 $Y=0.515 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_M1020_g N_VGND_c_660_n 0.00434272f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A_27_74#_M1021_g N_VGND_c_660_n 0.00434272f $X=5.195 $Y=0.74 $X2=0
+ $Y2=0
cc_313 N_A_27_74#_M1000_g N_VGND_c_663_n 0.0075754f $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A_27_74#_M1002_g N_VGND_c_663_n 0.0075754f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A_27_74#_M1006_g N_VGND_c_663_n 0.00820718f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A_27_74#_M1012_g N_VGND_c_663_n 0.00821294f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A_27_74#_M1016_g N_VGND_c_663_n 0.00821294f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_27_74#_M1017_g N_VGND_c_663_n 0.00821294f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A_27_74#_M1020_g N_VGND_c_663_n 0.00821344f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_27_74#_M1021_g N_VGND_c_663_n 0.00823984f $X=5.195 $Y=0.74 $X2=0
+ $Y2=0
cc_321 N_A_27_74#_c_178_n N_VGND_c_663_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_322 N_A_27_74#_c_181_n N_VGND_c_663_n 0.0062048f $X=1.185 $Y=0.515 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_403_n N_X_c_502_n 0.0256025f $X=1.635 $Y=2.455 $X2=0 $Y2=0
cc_324 N_VPWR_c_404_n N_X_c_502_n 0.0563525f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_325 N_VPWR_c_410_n N_X_c_502_n 0.0145938f $X=2.5 $Y=3.33 $X2=0 $Y2=0
cc_326 N_VPWR_c_401_n N_X_c_502_n 0.0120466f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_M1008_s N_X_c_503_n 0.00275645f $X=2.435 $Y=1.84 $X2=0 $Y2=0
cc_328 N_VPWR_c_404_n N_X_c_503_n 0.0184684f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_329 N_VPWR_c_404_n N_X_c_505_n 0.0322767f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_330 N_VPWR_c_405_n N_X_c_505_n 0.0563525f $X=3.535 $Y=2.305 $X2=0 $Y2=0
cc_331 N_VPWR_c_411_n N_X_c_505_n 0.014552f $X=3.45 $Y=3.33 $X2=0 $Y2=0
cc_332 N_VPWR_c_401_n N_X_c_505_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_333 N_VPWR_M1010_s N_X_c_506_n 0.00275645f $X=3.385 $Y=1.84 $X2=0 $Y2=0
cc_334 N_VPWR_c_405_n N_X_c_506_n 0.0184684f $X=3.535 $Y=2.305 $X2=0 $Y2=0
cc_335 N_VPWR_c_405_n N_X_c_507_n 0.0322767f $X=3.535 $Y=2.305 $X2=0 $Y2=0
cc_336 N_VPWR_c_406_n N_X_c_507_n 0.0563525f $X=4.485 $Y=2.305 $X2=0 $Y2=0
cc_337 N_VPWR_c_412_n N_X_c_507_n 0.014552f $X=4.4 $Y=3.33 $X2=0 $Y2=0
cc_338 N_VPWR_c_401_n N_X_c_507_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_339 N_VPWR_M1013_s N_X_c_508_n 0.002597f $X=4.335 $Y=1.84 $X2=0 $Y2=0
cc_340 N_VPWR_c_406_n N_X_c_508_n 0.017248f $X=4.485 $Y=2.305 $X2=0 $Y2=0
cc_341 N_VPWR_c_408_n X 0.0109193f $X=5.435 $Y=1.985 $X2=0 $Y2=0
cc_342 N_VPWR_c_406_n X 0.0336582f $X=4.485 $Y=2.305 $X2=0 $Y2=0
cc_343 N_VPWR_c_408_n X 0.0691255f $X=5.435 $Y=1.985 $X2=0 $Y2=0
cc_344 N_VPWR_c_413_n X 0.014802f $X=5.35 $Y=3.33 $X2=0 $Y2=0
cc_345 N_VPWR_c_401_n X 0.0122072f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_346 N_X_c_491_n N_VGND_M1002_s 0.00250873f $X=2.81 $Y=1.045 $X2=0 $Y2=0
cc_347 N_X_c_494_n N_VGND_M1012_s 0.00374767f $X=3.81 $Y=1.045 $X2=0 $Y2=0
cc_348 N_X_c_496_n N_VGND_M1017_s 0.00374767f $X=4.81 $Y=1.045 $X2=0 $Y2=0
cc_349 N_X_c_490_n N_VGND_c_646_n 0.0182488f $X=2.045 $Y=0.515 $X2=0 $Y2=0
cc_350 N_X_c_490_n N_VGND_c_647_n 0.0164567f $X=2.045 $Y=0.515 $X2=0 $Y2=0
cc_351 N_X_c_491_n N_VGND_c_647_n 0.0209867f $X=2.81 $Y=1.045 $X2=0 $Y2=0
cc_352 N_X_c_493_n N_VGND_c_647_n 0.0173003f $X=2.975 $Y=0.515 $X2=0 $Y2=0
cc_353 N_X_c_493_n N_VGND_c_648_n 0.0173003f $X=2.975 $Y=0.515 $X2=0 $Y2=0
cc_354 N_X_c_494_n N_VGND_c_648_n 0.0248957f $X=3.81 $Y=1.045 $X2=0 $Y2=0
cc_355 N_X_c_495_n N_VGND_c_648_n 0.0173003f $X=3.975 $Y=0.515 $X2=0 $Y2=0
cc_356 N_X_c_495_n N_VGND_c_649_n 0.0173003f $X=3.975 $Y=0.515 $X2=0 $Y2=0
cc_357 N_X_c_496_n N_VGND_c_649_n 0.0248957f $X=4.81 $Y=1.045 $X2=0 $Y2=0
cc_358 N_X_c_497_n N_VGND_c_649_n 0.0173384f $X=4.975 $Y=0.515 $X2=0 $Y2=0
cc_359 N_X_c_497_n N_VGND_c_651_n 0.0236943f $X=4.975 $Y=0.515 $X2=0 $Y2=0
cc_360 N_X_c_501_n N_VGND_c_651_n 0.00795492f $X=4.977 $Y=1.045 $X2=0 $Y2=0
cc_361 N_X_c_490_n N_VGND_c_652_n 0.00749631f $X=2.045 $Y=0.515 $X2=0 $Y2=0
cc_362 N_X_c_493_n N_VGND_c_654_n 0.0144922f $X=2.975 $Y=0.515 $X2=0 $Y2=0
cc_363 N_X_c_495_n N_VGND_c_656_n 0.0144922f $X=3.975 $Y=0.515 $X2=0 $Y2=0
cc_364 N_X_c_497_n N_VGND_c_660_n 0.0147153f $X=4.975 $Y=0.515 $X2=0 $Y2=0
cc_365 N_X_c_490_n N_VGND_c_663_n 0.0062048f $X=2.045 $Y=0.515 $X2=0 $Y2=0
cc_366 N_X_c_493_n N_VGND_c_663_n 0.0118826f $X=2.975 $Y=0.515 $X2=0 $Y2=0
cc_367 N_X_c_495_n N_VGND_c_663_n 0.0118826f $X=3.975 $Y=0.515 $X2=0 $Y2=0
cc_368 N_X_c_497_n N_VGND_c_663_n 0.0120673f $X=4.975 $Y=0.515 $X2=0 $Y2=0
