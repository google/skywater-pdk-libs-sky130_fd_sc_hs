* File: sky130_fd_sc_hs__clkdlyinv3sd2_1.pxi.spice
* Created: Tue Sep  1 19:58:05 2020
* 
x_PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A N_A_M1003_g N_A_c_51_n N_A_c_55_n
+ N_A_M1000_g A A N_A_c_53_n PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A
x_PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A_28_74# N_A_28_74#_M1003_s
+ N_A_28_74#_M1000_s N_A_28_74#_M1004_g N_A_28_74#_M1002_g N_A_28_74#_c_88_n
+ N_A_28_74#_c_94_n N_A_28_74#_c_95_n N_A_28_74#_c_104_n N_A_28_74#_c_89_n
+ N_A_28_74#_c_90_n N_A_28_74#_c_91_n N_A_28_74#_c_92_n
+ PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A_28_74#
x_PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A_288_74# N_A_288_74#_M1002_d
+ N_A_288_74#_M1004_d N_A_288_74#_M1005_g N_A_288_74#_c_150_n
+ N_A_288_74#_M1001_g N_A_288_74#_c_151_n N_A_288_74#_c_152_n
+ N_A_288_74#_c_153_n N_A_288_74#_c_157_n N_A_288_74#_c_154_n
+ PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A_288_74#
x_PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_s
+ N_VPWR_c_191_n N_VPWR_c_192_n VPWR N_VPWR_c_193_n N_VPWR_c_194_n
+ N_VPWR_c_195_n N_VPWR_c_190_n N_VPWR_c_197_n N_VPWR_c_198_n VPWR
+ PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%VPWR
x_PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%Y N_Y_M1005_d N_Y_M1001_d Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%Y
x_PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%VGND N_VGND_M1003_d N_VGND_M1005_s
+ N_VGND_c_239_n N_VGND_c_240_n VGND N_VGND_c_241_n N_VGND_c_242_n
+ N_VGND_c_243_n N_VGND_c_244_n N_VGND_c_245_n N_VGND_c_246_n VGND
+ PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%VGND
cc_1 VNB N_A_M1003_g 0.0470899f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.58
cc_2 VNB N_A_c_51_n 0.00890285f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.675
cc_3 VNB A 0.0265853f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_53_n 0.035867f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_5 VNB N_A_28_74#_M1002_g 0.0379702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_28_74#_c_88_n 0.0226356f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_7 VNB N_A_28_74#_c_89_n 0.0206633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_28_74#_c_90_n 0.0121635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_28_74#_c_91_n 0.00140945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_28_74#_c_92_n 0.0620251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_288_74#_M1005_g 0.0498775f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_12 VNB N_A_288_74#_c_150_n 0.0405564f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_A_288_74#_c_151_n 0.0216199f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_14 VNB N_A_288_74#_c_152_n 9.82213e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_288_74#_c_153_n 0.0209993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_288_74#_c_154_n 0.00614997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_190_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB Y 0.0204118f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_19 VNB Y 0.0485447f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_20 VNB N_VGND_c_239_n 0.00987431f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_21 VNB N_VGND_c_240_n 0.0107907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_241_n 0.0180717f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_23 VNB N_VGND_c_242_n 0.0303216f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.355
cc_24 VNB N_VGND_c_243_n 0.0187864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_244_n 0.191415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_245_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_246_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A_c_51_n 8.9669e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.675
cc_29 VPB N_A_c_55_n 0.0286196f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_30 VPB A 0.0106824f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_31 VPB N_A_28_74#_M1004_g 0.0362801f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_32 VPB N_A_28_74#_c_94_n 0.0079884f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.295
cc_33 VPB N_A_28_74#_c_95_n 0.0205617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_28_74#_c_91_n 0.00240258f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_28_74#_c_92_n 0.0135638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A_288_74#_c_150_n 0.0275939f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_37 VPB N_A_288_74#_c_152_n 0.0144837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_288_74#_c_157_n 0.00262425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_191_n 0.0101831f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_40 VPB N_VPWR_c_192_n 0.0174261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_193_n 0.018958f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.295
cc_42 VPB N_VPWR_c_194_n 0.0305232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_195_n 0.0182851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_190_n 0.0738836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_197_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_198_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB Y 0.00855207f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_48 VPB Y 0.0118233f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_49 VPB Y 0.0486918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 A N_A_28_74#_M1000_s 0.00256075f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_51 N_A_c_55_n N_A_28_74#_M1004_g 0.0140815f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_52 A N_A_28_74#_M1004_g 4.27742e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_53 N_A_M1003_g N_A_28_74#_M1002_g 0.00808739f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_54 N_A_M1003_g N_A_28_74#_c_88_n 0.0127782f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_55 A N_A_28_74#_c_94_n 0.0237727f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A_c_55_n N_A_28_74#_c_104_n 0.0144812f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_57 A N_A_28_74#_c_104_n 0.0197054f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_58 N_A_c_53_n N_A_28_74#_c_104_n 6.00585e-19 $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_59 N_A_M1003_g N_A_28_74#_c_89_n 0.0120856f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_60 A N_A_28_74#_c_89_n 0.0251751f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_A_c_53_n N_A_28_74#_c_89_n 0.00146806f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_62 N_A_M1003_g N_A_28_74#_c_90_n 0.00415005f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_63 A N_A_28_74#_c_90_n 0.0289843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A_M1003_g N_A_28_74#_c_91_n 0.0025292f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_65 N_A_c_51_n N_A_28_74#_c_91_n 2.04558e-19 $X=0.495 $Y=1.675 $X2=0 $Y2=0
cc_66 N_A_c_55_n N_A_28_74#_c_91_n 0.00383622f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_67 A N_A_28_74#_c_91_n 0.0416089f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_c_53_n N_A_28_74#_c_91_n 0.00110303f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_69 N_A_M1003_g N_A_28_74#_c_92_n 0.0021171f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_70 N_A_c_51_n N_A_28_74#_c_92_n 0.00643472f $X=0.495 $Y=1.675 $X2=0 $Y2=0
cc_71 A N_A_28_74#_c_92_n 0.00306446f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_c_53_n N_A_28_74#_c_92_n 0.0208886f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_73 A N_VPWR_M1000_d 0.00135779f $X=0.155 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_74 N_A_c_55_n N_VPWR_c_191_n 0.00426168f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A_c_55_n N_VPWR_c_193_n 0.00461464f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_c_55_n N_VPWR_c_190_n 0.00913361f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_VGND_c_239_n 0.00293875f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_78 N_A_M1003_g N_VGND_c_241_n 0.00456766f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_79 N_A_M1003_g N_VGND_c_244_n 0.00456437f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_80 N_A_28_74#_c_92_n N_A_288_74#_c_150_n 0.00356236f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_81 N_A_28_74#_M1002_g N_A_288_74#_c_151_n 0.0110261f $X=1.35 $Y=0.58 $X2=0
+ $Y2=0
cc_82 N_A_28_74#_c_89_n N_A_288_74#_c_151_n 0.0164122f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_83 N_A_28_74#_c_91_n N_A_288_74#_c_151_n 0.0211406f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_84 N_A_28_74#_c_92_n N_A_288_74#_c_151_n 0.0047987f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_85 N_A_28_74#_c_91_n N_A_288_74#_c_152_n 0.0285613f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_86 N_A_28_74#_c_92_n N_A_288_74#_c_152_n 0.00885412f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_87 N_A_28_74#_M1004_g N_A_288_74#_c_157_n 0.00707225f $X=1.32 $Y=2.46 $X2=0
+ $Y2=0
cc_88 N_A_28_74#_c_91_n N_A_288_74#_c_154_n 0.0278254f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_89 N_A_28_74#_c_92_n N_A_288_74#_c_154_n 0.00523717f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_90 N_A_28_74#_c_104_n N_VPWR_M1000_d 0.0249816f $X=0.975 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_28_74#_c_91_n N_VPWR_M1000_d 0.0012063f $X=1.14 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_28_74#_M1004_g N_VPWR_c_191_n 0.0104916f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_93 N_A_28_74#_c_104_n N_VPWR_c_191_n 0.0220956f $X=0.975 $Y=2.117 $X2=0 $Y2=0
cc_94 N_A_28_74#_M1004_g N_VPWR_c_192_n 0.0044498f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_95 N_A_28_74#_c_95_n N_VPWR_c_193_n 0.00593336f $X=0.265 $Y=2.56 $X2=0 $Y2=0
cc_96 N_A_28_74#_M1004_g N_VPWR_c_194_n 0.00738282f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_97 N_A_28_74#_M1004_g N_VPWR_c_190_n 0.014148f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_98 N_A_28_74#_c_95_n N_VPWR_c_190_n 0.00940928f $X=0.265 $Y=2.56 $X2=0 $Y2=0
cc_99 N_A_28_74#_M1002_g N_VGND_c_239_n 0.00513169f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_100 N_A_28_74#_c_88_n N_VGND_c_239_n 0.0151665f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_101 N_A_28_74#_c_89_n N_VGND_c_239_n 0.0255952f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_102 N_A_28_74#_M1002_g N_VGND_c_240_n 0.00247044f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_103 N_A_28_74#_c_88_n N_VGND_c_241_n 0.0170785f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_104 N_A_28_74#_M1002_g N_VGND_c_242_n 0.00553757f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_105 N_A_28_74#_M1002_g N_VGND_c_244_n 0.00962875f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_106 N_A_28_74#_c_88_n N_VGND_c_244_n 0.0118627f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_107 N_A_28_74#_c_89_n N_VGND_c_244_n 0.0213669f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_108 N_A_288_74#_c_157_n N_VPWR_c_191_n 0.00825858f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_109 N_A_288_74#_c_150_n N_VPWR_c_192_n 0.0193941f $X=2.325 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_288_74#_c_152_n N_VPWR_c_192_n 0.0761011f $X=1.58 $Y=2.105 $X2=0
+ $Y2=0
cc_111 N_A_288_74#_c_153_n N_VPWR_c_192_n 0.0176738f $X=2.275 $Y=1.46 $X2=0
+ $Y2=0
cc_112 N_A_288_74#_c_157_n N_VPWR_c_194_n 0.00976575f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_113 N_A_288_74#_c_150_n N_VPWR_c_195_n 0.00413917f $X=2.325 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_288_74#_c_150_n N_VPWR_c_190_n 0.00821375f $X=2.325 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_288_74#_c_157_n N_VPWR_c_190_n 0.0112865f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_116 N_A_288_74#_M1005_g Y 8.21909e-19 $X=2.315 $Y=0.58 $X2=0 $Y2=0
cc_117 N_A_288_74#_M1005_g Y 0.0195788f $X=2.315 $Y=0.58 $X2=0 $Y2=0
cc_118 N_A_288_74#_c_150_n Y 0.0155759f $X=2.325 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_288_74#_c_153_n Y 0.0270738f $X=2.275 $Y=1.46 $X2=0 $Y2=0
cc_120 N_A_288_74#_c_150_n Y 0.00443902f $X=2.325 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_288_74#_c_151_n N_VGND_c_239_n 0.00689121f $X=1.58 $Y=0.58 $X2=0
+ $Y2=0
cc_122 N_A_288_74#_M1005_g N_VGND_c_240_n 0.0132522f $X=2.315 $Y=0.58 $X2=0
+ $Y2=0
cc_123 N_A_288_74#_c_150_n N_VGND_c_240_n 0.00210741f $X=2.325 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_288_74#_c_151_n N_VGND_c_240_n 0.0307431f $X=1.58 $Y=0.58 $X2=0 $Y2=0
cc_125 N_A_288_74#_c_153_n N_VGND_c_240_n 0.0105553f $X=2.275 $Y=1.46 $X2=0
+ $Y2=0
cc_126 N_A_288_74#_c_151_n N_VGND_c_242_n 0.0132196f $X=1.58 $Y=0.58 $X2=0 $Y2=0
cc_127 N_A_288_74#_M1005_g N_VGND_c_243_n 0.00383152f $X=2.315 $Y=0.58 $X2=0
+ $Y2=0
cc_128 N_A_288_74#_M1005_g N_VGND_c_244_n 0.00761414f $X=2.315 $Y=0.58 $X2=0
+ $Y2=0
cc_129 N_A_288_74#_c_151_n N_VGND_c_244_n 0.00920999f $X=1.58 $Y=0.58 $X2=0
+ $Y2=0
cc_130 N_VPWR_c_192_n Y 0.0476994f $X=2.1 $Y=1.985 $X2=0 $Y2=0
cc_131 N_VPWR_c_195_n Y 0.0234396f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_132 N_VPWR_c_190_n Y 0.0138183f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_133 Y N_VGND_c_240_n 0.0154115f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_134 Y N_VGND_c_243_n 0.0155069f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_135 Y N_VGND_c_244_n 0.013122f $X=2.555 $Y=0.47 $X2=0 $Y2=0
