* File: sky130_fd_sc_hs__o41ai_2.spice
* Created: Tue Sep  1 20:19:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o41ai_2.pex.spice"
.subckt sky130_fd_sc_hs__o41ai_2  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_A_132_74#_M1008_d N_B1_M1008_g N_Y_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75004.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_132_74#_M1018_d N_B1_M1018_g N_Y_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75004.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_132_74#_M1018_d N_A4_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1006 N_A_132_74#_M1006_d N_A4_M1006_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12765 AS=0.1295 PD=1.085 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A3_M1011_g N_A_132_74#_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.12765 PD=1.025 PS=1.085 NRD=0.804 NRS=10.536 M=1 R=4.93333
+ SA=75002.1 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1011_d N_A3_M1012_g N_A_132_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.1147 PD=1.025 PS=1.05 NRD=0 NRS=2.424 M=1 R=4.93333 SA=75002.6
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1013 N_A_132_74#_M1012_s N_A2_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1554 PD=1.05 PS=1.16 NRD=2.424 NRS=11.34 M=1 R=4.93333 SA=75003
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1017 N_A_132_74#_M1017_d N_A2_M1017_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_132_74#_M1017_d N_A1_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1016 N_A_132_74#_M1016_d N_A1_M1016_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1295 PD=2.19 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.5
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1001_d N_B1_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3136 PD=1.42 PS=2.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75000.2 A=0.168 P=2.54 MULT=1
MM1003 N_A_314_368#_M1003_d N_A4_M1003_g N_Y_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3136 AS=0.168 PD=2.8 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1019 N_A_314_368#_M1019_d N_A4_M1019_g N_Y_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2436 AS=0.168 PD=1.555 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1007 N_A_607_368#_M1007_d N_A3_M1007_g N_A_314_368#_M1019_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.2436 PD=1.42 PS=1.555 NRD=1.7533 NRS=25.4918 M=1
+ R=7.46667 SA=75001.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_A_607_368#_M1007_d N_A3_M1009_g N_A_314_368#_M1009_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3136 PD=1.42 PS=2.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_607_368#_M1000_d N_A2_M1000_g N_A_807_368#_M1000_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1004 N_A_607_368#_M1000_d N_A2_M1004_g N_A_807_368#_M1004_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_807_368#_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1010_d N_A1_M1014_g N_A_807_368#_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3132 P=16.96
c_111 VPB 0 1.5035e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__o41ai_2.pxi.spice"
*
.ends
*
*
