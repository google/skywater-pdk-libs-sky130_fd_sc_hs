* File: sky130_fd_sc_hs__sdfrtp_1.pxi.spice
* Created: Tue Sep  1 20:22:38 2020
* 
x_PM_SKY130_FD_SC_HS__SDFRTP_1%SCE N_SCE_c_298_n N_SCE_M1037_g N_SCE_c_299_n
+ N_SCE_M1023_g N_SCE_c_300_n N_SCE_c_301_n N_SCE_M1020_g N_SCE_M1030_g
+ N_SCE_c_293_n N_SCE_c_294_n N_SCE_c_295_n SCE SCE SCE N_SCE_c_296_n
+ N_SCE_c_297_n SCE N_SCE_c_305_n PM_SKY130_FD_SC_HS__SDFRTP_1%SCE
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_27_88# N_A_27_88#_M1037_s N_A_27_88#_M1023_s
+ N_A_27_88#_c_378_n N_A_27_88#_M1012_g N_A_27_88#_c_385_n N_A_27_88#_M1024_g
+ N_A_27_88#_c_379_n N_A_27_88#_c_380_n N_A_27_88#_c_387_n N_A_27_88#_c_381_n
+ N_A_27_88#_c_388_n N_A_27_88#_c_389_n N_A_27_88#_c_390_n N_A_27_88#_c_382_n
+ N_A_27_88#_c_391_n N_A_27_88#_c_383_n N_A_27_88#_c_384_n N_A_27_88#_c_392_n
+ PM_SKY130_FD_SC_HS__SDFRTP_1%A_27_88#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%D N_D_c_468_n N_D_M1036_g N_D_c_462_n N_D_c_463_n
+ N_D_M1013_g N_D_c_470_n N_D_c_464_n D N_D_c_465_n N_D_c_466_n N_D_c_467_n
+ PM_SKY130_FD_SC_HS__SDFRTP_1%D
x_PM_SKY130_FD_SC_HS__SDFRTP_1%SCD N_SCD_c_520_n N_SCD_M1006_g N_SCD_M1021_g
+ N_SCD_c_517_n SCD SCD N_SCD_c_519_n PM_SKY130_FD_SC_HS__SDFRTP_1%SCD
x_PM_SKY130_FD_SC_HS__SDFRTP_1%RESET_B N_RESET_B_c_568_n N_RESET_B_M1039_g
+ N_RESET_B_M1016_g N_RESET_B_c_561_n N_RESET_B_M1019_g N_RESET_B_c_562_n
+ N_RESET_B_c_563_n N_RESET_B_c_564_n N_RESET_B_c_571_n N_RESET_B_M1034_g
+ N_RESET_B_M1038_g N_RESET_B_c_566_n N_RESET_B_c_573_n N_RESET_B_c_574_n
+ N_RESET_B_M1015_g N_RESET_B_c_567_n N_RESET_B_c_575_n N_RESET_B_c_576_n
+ N_RESET_B_c_577_n N_RESET_B_c_578_n N_RESET_B_c_579_n RESET_B
+ N_RESET_B_c_581_n N_RESET_B_c_582_n N_RESET_B_c_583_n N_RESET_B_c_584_n
+ N_RESET_B_c_585_n PM_SKY130_FD_SC_HS__SDFRTP_1%RESET_B
x_PM_SKY130_FD_SC_HS__SDFRTP_1%CLK N_CLK_c_772_n N_CLK_M1022_g N_CLK_M1008_g
+ N_CLK_c_774_n N_CLK_c_785_n CLK N_CLK_c_775_n PM_SKY130_FD_SC_HS__SDFRTP_1%CLK
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_1034_368# N_A_1034_368#_M1003_d
+ N_A_1034_368#_M1029_d N_A_1034_368#_c_845_n N_A_1034_368#_c_846_n
+ N_A_1034_368#_M1026_g N_A_1034_368#_c_824_n N_A_1034_368#_M1000_g
+ N_A_1034_368#_c_826_n N_A_1034_368#_M1010_g N_A_1034_368#_c_827_n
+ N_A_1034_368#_c_848_n N_A_1034_368#_M1025_g N_A_1034_368#_c_828_n
+ N_A_1034_368#_c_829_n N_A_1034_368#_c_830_n N_A_1034_368#_c_831_n
+ N_A_1034_368#_c_832_n N_A_1034_368#_c_833_n N_A_1034_368#_c_834_n
+ N_A_1034_368#_c_835_n N_A_1034_368#_c_872_p N_A_1034_368#_c_862_n
+ N_A_1034_368#_c_836_n N_A_1034_368#_c_837_n N_A_1034_368#_c_838_n
+ N_A_1034_368#_c_839_n N_A_1034_368#_c_961_p N_A_1034_368#_c_852_n
+ N_A_1034_368#_c_840_n N_A_1034_368#_c_841_n N_A_1034_368#_c_842_n
+ N_A_1034_368#_c_843_n N_A_1034_368#_c_844_n
+ PM_SKY130_FD_SC_HS__SDFRTP_1%A_1034_368#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_1367_92# N_A_1367_92#_M1033_d
+ N_A_1367_92#_M1001_d N_A_1367_92#_M1027_g N_A_1367_92#_c_1044_n
+ N_A_1367_92#_c_1045_n N_A_1367_92#_M1002_g N_A_1367_92#_c_1038_n
+ N_A_1367_92#_c_1039_n N_A_1367_92#_c_1040_n N_A_1367_92#_c_1041_n
+ N_A_1367_92#_c_1048_n N_A_1367_92#_c_1049_n N_A_1367_92#_c_1042_n
+ N_A_1367_92#_c_1043_n PM_SKY130_FD_SC_HS__SDFRTP_1%A_1367_92#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_1233_118# N_A_1233_118#_M1009_d
+ N_A_1233_118#_M1026_d N_A_1233_118#_M1034_d N_A_1233_118#_M1033_g
+ N_A_1233_118#_c_1147_n N_A_1233_118#_c_1156_n N_A_1233_118#_M1001_g
+ N_A_1233_118#_c_1157_n N_A_1233_118#_c_1148_n N_A_1233_118#_c_1149_n
+ N_A_1233_118#_c_1168_n N_A_1233_118#_c_1150_n N_A_1233_118#_c_1151_n
+ N_A_1233_118#_c_1152_n N_A_1233_118#_c_1153_n N_A_1233_118#_c_1154_n
+ N_A_1233_118#_c_1161_n PM_SKY130_FD_SC_HS__SDFRTP_1%A_1233_118#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_855_368# N_A_855_368#_M1008_s
+ N_A_855_368#_M1022_s N_A_855_368#_c_1280_n N_A_855_368#_M1029_g
+ N_A_855_368#_c_1281_n N_A_855_368#_M1003_g N_A_855_368#_c_1282_n
+ N_A_855_368#_c_1283_n N_A_855_368#_c_1284_n N_A_855_368#_c_1298_n
+ N_A_855_368#_c_1299_n N_A_855_368#_M1009_g N_A_855_368#_c_1300_n
+ N_A_855_368#_c_1301_n N_A_855_368#_c_1302_n N_A_855_368#_M1032_g
+ N_A_855_368#_c_1303_n N_A_855_368#_c_1304_n N_A_855_368#_c_1305_n
+ N_A_855_368#_M1004_g N_A_855_368#_c_1286_n N_A_855_368#_c_1287_n
+ N_A_855_368#_c_1288_n N_A_855_368#_M1007_g N_A_855_368#_c_1290_n
+ N_A_855_368#_c_1309_n N_A_855_368#_c_1291_n N_A_855_368#_c_1292_n
+ N_A_855_368#_c_1336_n N_A_855_368#_c_1322_n N_A_855_368#_c_1310_n
+ N_A_855_368#_c_1293_n N_A_855_368#_c_1294_n N_A_855_368#_c_1312_n
+ N_A_855_368#_c_1295_n PM_SKY130_FD_SC_HS__SDFRTP_1%A_855_368#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_1997_272# N_A_1997_272#_M1028_d
+ N_A_1997_272#_M1015_d N_A_1997_272#_M1005_g N_A_1997_272#_c_1483_n
+ N_A_1997_272#_c_1494_n N_A_1997_272#_c_1495_n N_A_1997_272#_M1014_g
+ N_A_1997_272#_c_1484_n N_A_1997_272#_c_1485_n N_A_1997_272#_c_1486_n
+ N_A_1997_272#_c_1487_n N_A_1997_272#_c_1488_n N_A_1997_272#_c_1489_n
+ N_A_1997_272#_c_1490_n N_A_1997_272#_c_1496_n N_A_1997_272#_c_1491_n
+ N_A_1997_272#_c_1492_n PM_SKY130_FD_SC_HS__SDFRTP_1%A_1997_272#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_1745_74# N_A_1745_74#_M1010_d
+ N_A_1745_74#_M1004_d N_A_1745_74#_M1028_g N_A_1745_74#_c_1600_n
+ N_A_1745_74#_c_1611_n N_A_1745_74#_c_1612_n N_A_1745_74#_M1018_g
+ N_A_1745_74#_c_1601_n N_A_1745_74#_c_1602_n N_A_1745_74#_c_1613_n
+ N_A_1745_74#_c_1614_n N_A_1745_74#_M1017_g N_A_1745_74#_M1031_g
+ N_A_1745_74#_c_1615_n N_A_1745_74#_c_1616_n N_A_1745_74#_c_1604_n
+ N_A_1745_74#_c_1605_n N_A_1745_74#_c_1618_n N_A_1745_74#_c_1619_n
+ N_A_1745_74#_c_1620_n N_A_1745_74#_c_1606_n N_A_1745_74#_c_1607_n
+ N_A_1745_74#_c_1608_n N_A_1745_74#_c_1609_n
+ PM_SKY130_FD_SC_HS__SDFRTP_1%A_1745_74#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_2399_424# N_A_2399_424#_M1031_d
+ N_A_2399_424#_M1017_d N_A_2399_424#_c_1771_n N_A_2399_424#_M1035_g
+ N_A_2399_424#_M1011_g N_A_2399_424#_c_1767_n N_A_2399_424#_c_1773_n
+ N_A_2399_424#_c_1768_n N_A_2399_424#_c_1793_p N_A_2399_424#_c_1769_n
+ N_A_2399_424#_c_1770_n PM_SKY130_FD_SC_HS__SDFRTP_1%A_2399_424#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%VPWR N_VPWR_M1023_d N_VPWR_M1006_d N_VPWR_M1022_d
+ N_VPWR_M1002_d N_VPWR_M1001_s N_VPWR_M1014_d N_VPWR_M1018_d N_VPWR_M1035_s
+ N_VPWR_c_1814_n N_VPWR_c_1815_n N_VPWR_c_1816_n N_VPWR_c_1817_n
+ N_VPWR_c_1818_n N_VPWR_c_1819_n N_VPWR_c_1820_n N_VPWR_c_1821_n
+ N_VPWR_c_1822_n N_VPWR_c_1823_n N_VPWR_c_1824_n N_VPWR_c_1825_n
+ N_VPWR_c_1826_n N_VPWR_c_1827_n N_VPWR_c_1828_n VPWR N_VPWR_c_1829_n
+ N_VPWR_c_1830_n N_VPWR_c_1831_n N_VPWR_c_1832_n N_VPWR_c_1833_n
+ N_VPWR_c_1813_n N_VPWR_c_1835_n N_VPWR_c_1836_n N_VPWR_c_1837_n
+ N_VPWR_c_1838_n N_VPWR_c_1839_n PM_SKY130_FD_SC_HS__SDFRTP_1%VPWR
x_PM_SKY130_FD_SC_HS__SDFRTP_1%A_300_464# N_A_300_464#_M1013_d
+ N_A_300_464#_M1009_s N_A_300_464#_M1036_d N_A_300_464#_M1039_d
+ N_A_300_464#_M1026_s N_A_300_464#_c_1982_n N_A_300_464#_c_2001_n
+ N_A_300_464#_c_1975_n N_A_300_464#_c_1976_n N_A_300_464#_c_1984_n
+ N_A_300_464#_c_1985_n N_A_300_464#_c_1977_n N_A_300_464#_c_1986_n
+ N_A_300_464#_c_1978_n N_A_300_464#_c_1979_n N_A_300_464#_c_1987_n
+ N_A_300_464#_c_1988_n N_A_300_464#_c_1980_n N_A_300_464#_c_1990_n
+ N_A_300_464#_c_1981_n N_A_300_464#_c_1991_n
+ PM_SKY130_FD_SC_HS__SDFRTP_1%A_300_464#
x_PM_SKY130_FD_SC_HS__SDFRTP_1%Q N_Q_M1011_d N_Q_M1035_d Q Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_HS__SDFRTP_1%Q
x_PM_SKY130_FD_SC_HS__SDFRTP_1%VGND N_VGND_M1037_d N_VGND_M1016_d N_VGND_M1008_d
+ N_VGND_M1019_d N_VGND_M1005_d N_VGND_M1031_s N_VGND_M1011_s N_VGND_c_2147_n
+ N_VGND_c_2148_n N_VGND_c_2149_n N_VGND_c_2150_n N_VGND_c_2151_n
+ N_VGND_c_2152_n N_VGND_c_2153_n N_VGND_c_2154_n N_VGND_c_2155_n
+ N_VGND_c_2156_n VGND N_VGND_c_2157_n N_VGND_c_2158_n N_VGND_c_2159_n
+ N_VGND_c_2160_n N_VGND_c_2161_n N_VGND_c_2162_n N_VGND_c_2163_n
+ N_VGND_c_2164_n N_VGND_c_2165_n N_VGND_c_2166_n N_VGND_c_2167_n
+ N_VGND_c_2168_n PM_SKY130_FD_SC_HS__SDFRTP_1%VGND
x_PM_SKY130_FD_SC_HS__SDFRTP_1%noxref_24 N_noxref_24_M1012_s N_noxref_24_M1021_d
+ N_noxref_24_c_2273_n N_noxref_24_c_2274_n
+ PM_SKY130_FD_SC_HS__SDFRTP_1%noxref_24
cc_1 VNB N_SCE_M1037_g 0.062352f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_2 VNB N_SCE_M1030_g 0.0341303f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_3 VNB N_SCE_c_293_n 0.014614f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=1.575
cc_4 VNB N_SCE_c_294_n 0.00230215f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_5 VNB N_SCE_c_295_n 0.0345925f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_6 VNB N_SCE_c_296_n 0.0331371f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_7 VNB N_SCE_c_297_n 0.0110089f $X=-0.19 $Y=-0.245 $X2=1.623 $Y2=1.662
cc_8 VNB N_A_27_88#_c_378_n 0.0192577f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_9 VNB N_A_27_88#_c_379_n 0.0282802f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_10 VNB N_A_27_88#_c_380_n 0.0187337f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.575
cc_11 VNB N_A_27_88#_c_381_n 0.0167058f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.575
cc_12 VNB N_A_27_88#_c_382_n 0.0130086f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.67
cc_13 VNB N_A_27_88#_c_383_n 0.00840348f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_14 VNB N_A_27_88#_c_384_n 0.0522403f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_15 VNB N_D_c_462_n 0.00442527f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_16 VNB N_D_c_463_n 0.0153194f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_17 VNB N_D_c_464_n 0.021136f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.26
cc_18 VNB N_D_c_465_n 0.032448f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.575
cc_19 VNB N_D_c_466_n 0.00949867f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_20 VNB N_D_c_467_n 0.0161824f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_21 VNB N_SCD_M1021_g 0.0442872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCD_c_517_n 0.00430596f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.835
cc_23 VNB SCD 0.00223563f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.155
cc_24 VNB N_SCD_c_519_n 0.0171077f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_25 VNB N_RESET_B_M1016_g 0.0636082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_RESET_B_c_561_n 0.0166101f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_27 VNB N_RESET_B_c_562_n 0.0276292f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.155
cc_28 VNB N_RESET_B_c_563_n 0.0071197f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.245
cc_29 VNB N_RESET_B_c_564_n 0.0221058f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.64
cc_30 VNB N_RESET_B_M1038_g 0.0378564f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.575
cc_31 VNB N_RESET_B_c_566_n 0.0109809f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_32 VNB N_RESET_B_c_567_n 0.0164222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_CLK_c_772_n 0.0189694f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.835
cc_34 VNB N_CLK_M1008_g 0.0229621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_CLK_c_774_n 0.0596142f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_36 VNB N_CLK_c_775_n 0.0130134f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_37 VNB N_A_1034_368#_c_824_n 0.0100727f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.245
cc_38 VNB N_A_1034_368#_M1000_g 0.040778f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_39 VNB N_A_1034_368#_c_826_n 0.0161967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1034_368#_c_827_n 0.00792759f $X=-0.19 $Y=-0.245 $X2=2.56
+ $Y2=1.425
cc_41 VNB N_A_1034_368#_c_828_n 0.00792011f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=1.58
cc_42 VNB N_A_1034_368#_c_829_n 0.00211344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1034_368#_c_830_n 0.0441847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1034_368#_c_831_n 0.0046921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1034_368#_c_832_n 7.95232e-19 $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_46 VNB N_A_1034_368#_c_833_n 0.00175807f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_47 VNB N_A_1034_368#_c_834_n 0.00449285f $X=-0.19 $Y=-0.245 $X2=2.56
+ $Y2=1.425
cc_48 VNB N_A_1034_368#_c_835_n 8.10761e-19 $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.26
cc_49 VNB N_A_1034_368#_c_836_n 0.00889307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1034_368#_c_837_n 0.00245962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1034_368#_c_838_n 0.00270816f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.662
cc_52 VNB N_A_1034_368#_c_839_n 0.00419892f $X=-0.19 $Y=-0.245 $X2=1.609
+ $Y2=1.662
cc_53 VNB N_A_1034_368#_c_840_n 0.00503286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1034_368#_c_841_n 0.0363807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1034_368#_c_842_n 0.00354363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1034_368#_c_843_n 0.0117407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1034_368#_c_844_n 0.0259737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1367_92#_M1027_g 0.0336377f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_59 VNB N_A_1367_92#_c_1038_n 0.00388286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1367_92#_c_1039_n 0.0258247f $X=-0.19 $Y=-0.245 $X2=2.395
+ $Y2=1.575
cc_61 VNB N_A_1367_92#_c_1040_n 0.00326481f $X=-0.19 $Y=-0.245 $X2=2.56
+ $Y2=1.425
cc_62 VNB N_A_1367_92#_c_1041_n 4.68114e-19 $X=-0.19 $Y=-0.245 $X2=2.56
+ $Y2=1.425
cc_63 VNB N_A_1367_92#_c_1042_n 0.00364646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1367_92#_c_1043_n 0.00552017f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_65 VNB N_A_1233_118#_M1033_g 0.0261617f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.245
cc_66 VNB N_A_1233_118#_c_1147_n 0.0175736f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.64
cc_67 VNB N_A_1233_118#_c_1148_n 0.00391631f $X=-0.19 $Y=-0.245 $X2=2.56
+ $Y2=1.425
cc_68 VNB N_A_1233_118#_c_1149_n 0.00426083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1233_118#_c_1150_n 4.99311e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1233_118#_c_1151_n 0.00277903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1233_118#_c_1152_n 0.00602363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1233_118#_c_1153_n 0.0280028f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_73 VNB N_A_1233_118#_c_1154_n 0.00206355f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_74 VNB N_A_855_368#_c_1280_n 0.0334321f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.245
cc_75 VNB N_A_855_368#_c_1281_n 0.0179355f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.835
cc_76 VNB N_A_855_368#_c_1282_n 0.0127757f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.64
cc_77 VNB N_A_855_368#_c_1283_n 0.0142334f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_78 VNB N_A_855_368#_c_1284_n 0.0262621f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_79 VNB N_A_855_368#_M1009_g 0.0213501f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_80 VNB N_A_855_368#_c_1286_n 0.0179478f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_81 VNB N_A_855_368#_c_1287_n 0.00460795f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.67
cc_82 VNB N_A_855_368#_c_1288_n 0.0208108f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.26
cc_83 VNB N_A_855_368#_M1007_g 0.0235073f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.662
cc_84 VNB N_A_855_368#_c_1290_n 0.00856677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_855_368#_c_1291_n 0.0124432f $X=-0.19 $Y=-0.245 $X2=1.609
+ $Y2=1.662
cc_86 VNB N_A_855_368#_c_1292_n 0.00188799f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.662
cc_87 VNB N_A_855_368#_c_1293_n 0.00256459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_855_368#_c_1294_n 9.18582e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_855_368#_c_1295_n 0.00472377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1997_272#_M1005_g 0.0393068f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_91 VNB N_A_1997_272#_c_1483_n 0.0235946f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.155
cc_92 VNB N_A_1997_272#_c_1484_n 0.0152817f $X=-0.19 $Y=-0.245 $X2=2.65
+ $Y2=0.615
cc_93 VNB N_A_1997_272#_c_1485_n 0.0073172f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.575
cc_94 VNB N_A_1997_272#_c_1486_n 0.00658513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1997_272#_c_1487_n 0.00719764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1997_272#_c_1488_n 0.00239418f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_97 VNB N_A_1997_272#_c_1489_n 0.00890748f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=1.58
cc_98 VNB N_A_1997_272#_c_1490_n 0.00132368f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_99 VNB N_A_1997_272#_c_1491_n 4.91246e-19 $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_100 VNB N_A_1997_272#_c_1492_n 6.26987e-19 $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.67
cc_101 VNB N_A_1745_74#_M1028_g 0.0220606f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_102 VNB N_A_1745_74#_c_1600_n 0.0178723f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.245
cc_103 VNB N_A_1745_74#_c_1601_n 0.0372707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1745_74#_c_1602_n 0.0476514f $X=-0.19 $Y=-0.245 $X2=2.395
+ $Y2=1.575
cc_105 VNB N_A_1745_74#_M1031_g 0.0313727f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_106 VNB N_A_1745_74#_c_1604_n 0.0027518f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.67
cc_107 VNB N_A_1745_74#_c_1605_n 0.00220477f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_108 VNB N_A_1745_74#_c_1606_n 0.00284242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1745_74#_c_1607_n 0.00104193f $X=-0.19 $Y=-0.245 $X2=1.2
+ $Y2=1.662
cc_110 VNB N_A_1745_74#_c_1608_n 8.69032e-19 $X=-0.19 $Y=-0.245 $X2=1.609
+ $Y2=1.662
cc_111 VNB N_A_1745_74#_c_1609_n 0.0278597f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=1.665
cc_112 VNB N_A_2399_424#_M1011_g 0.0281108f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.245
cc_113 VNB N_A_2399_424#_c_1767_n 0.0900229f $X=-0.19 $Y=-0.245 $X2=2.65
+ $Y2=1.26
cc_114 VNB N_A_2399_424#_c_1768_n 0.016101f $X=-0.19 $Y=-0.245 $X2=2.56
+ $Y2=1.425
cc_115 VNB N_A_2399_424#_c_1769_n 8.47259e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2399_424#_c_1770_n 0.00458466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VPWR_c_1813_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_300_464#_c_1975_n 0.023632f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_119 VNB N_A_300_464#_c_1976_n 0.00514666f $X=-0.19 $Y=-0.245 $X2=2.56
+ $Y2=1.575
cc_120 VNB N_A_300_464#_c_1977_n 0.00283431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_300_464#_c_1978_n 0.0053476f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_122 VNB N_A_300_464#_c_1979_n 0.00160258f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_123 VNB N_A_300_464#_c_1980_n 0.00381868f $X=-0.19 $Y=-0.245 $X2=2.56
+ $Y2=1.26
cc_124 VNB N_A_300_464#_c_1981_n 0.00548504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB Q 0.0259999f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_126 VNB Q 0.00837931f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_127 VNB Q 0.027119f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_128 VNB N_VGND_c_2147_n 0.0181638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2148_n 0.00943648f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_130 VNB N_VGND_c_2149_n 0.00526449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2150_n 0.0100142f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_132 VNB N_VGND_c_2151_n 0.00854448f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.425
cc_133 VNB N_VGND_c_2152_n 0.0169646f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.662
cc_134 VNB N_VGND_c_2153_n 0.0690616f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.662
cc_135 VNB N_VGND_c_2154_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.662
cc_136 VNB N_VGND_c_2155_n 0.0226507f $X=-0.19 $Y=-0.245 $X2=1.609 $Y2=1.662
cc_137 VNB N_VGND_c_2156_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.662
cc_138 VNB N_VGND_c_2157_n 0.0177976f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.662
cc_139 VNB N_VGND_c_2158_n 0.057793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2159_n 0.0611983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2160_n 0.0297773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2161_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2162_n 0.0194697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2163_n 0.752337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2164_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2165_n 0.0148571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2166_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2167_n 0.00622769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2168_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_noxref_24_c_2273_n 0.01789f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_151 VNB N_noxref_24_c_2274_n 0.00667823f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.64
cc_152 VPB N_SCE_c_298_n 0.0195456f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.155
cc_153 VPB N_SCE_c_299_n 0.0273001f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_154 VPB N_SCE_c_300_n 0.0184657f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.155
cc_155 VPB N_SCE_c_301_n 0.02161f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_156 VPB N_SCE_c_294_n 0.00260547f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.425
cc_157 VPB N_SCE_c_296_n 0.0253807f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_158 VPB N_SCE_c_297_n 0.00455267f $X=-0.19 $Y=1.66 $X2=1.623 $Y2=1.662
cc_159 VPB N_SCE_c_305_n 0.00736556f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.662
cc_160 VPB N_A_27_88#_c_385_n 0.0422502f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_161 VPB N_A_27_88#_c_380_n 0.0161852f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.575
cc_162 VPB N_A_27_88#_c_387_n 0.0338402f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.425
cc_163 VPB N_A_27_88#_c_388_n 0.00369885f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_164 VPB N_A_27_88#_c_389_n 0.00550456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_27_88#_c_390_n 0.0465306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_27_88#_c_391_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.67
cc_167 VPB N_A_27_88#_c_392_n 0.0240446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_D_c_468_n 0.0213045f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.835
cc_169 VPB N_D_c_462_n 0.0250339f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.65
cc_170 VPB N_D_c_470_n 0.029832f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.155
cc_171 VPB N_SCD_c_520_n 0.0161432f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.835
cc_172 VPB N_SCD_c_517_n 0.051049f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.835
cc_173 VPB SCD 0.00172059f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.155
cc_174 VPB N_RESET_B_c_568_n 0.0424629f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.835
cc_175 VPB N_RESET_B_M1016_g 0.0129227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_RESET_B_c_564_n 0.010477f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_177 VPB N_RESET_B_c_571_n 0.0167021f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=1.26
cc_178 VPB N_RESET_B_c_566_n 0.00936563f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.425
cc_179 VPB N_RESET_B_c_573_n 0.0136009f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.575
cc_180 VPB N_RESET_B_c_574_n 0.0233932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_RESET_B_c_575_n 0.0234239f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.67
cc_182 VPB N_RESET_B_c_576_n 0.00161953f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_183 VPB N_RESET_B_c_577_n 0.0217281f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_184 VPB N_RESET_B_c_578_n 0.0020849f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_185 VPB N_RESET_B_c_579_n 0.00628945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB RESET_B 0.00299651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_RESET_B_c_581_n 0.0437469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_RESET_B_c_582_n 0.00233009f $X=-0.19 $Y=1.66 $X2=1.609 $Y2=1.662
cc_189 VPB N_RESET_B_c_583_n 0.0598827f $X=-0.19 $Y=1.66 $X2=1.694 $Y2=1.662
cc_190 VPB N_RESET_B_c_584_n 0.00324614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_RESET_B_c_585_n 0.0327579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_CLK_c_772_n 0.0297766f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.835
cc_193 VPB N_A_1034_368#_c_845_n 0.0159039f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_194 VPB N_A_1034_368#_c_846_n 0.0203624f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_195 VPB N_A_1034_368#_c_824_n 0.0136311f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_196 VPB N_A_1034_368#_c_848_n 0.0607238f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.425
cc_197 VPB N_A_1034_368#_c_832_n 0.0074594f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.67
cc_198 VPB N_A_1034_368#_c_833_n 0.00200713f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_199 VPB N_A_1034_368#_c_839_n 0.00116335f $X=-0.19 $Y=1.66 $X2=1.609
+ $Y2=1.662
cc_200 VPB N_A_1034_368#_c_852_n 0.00218598f $X=-0.19 $Y=1.66 $X2=1.694
+ $Y2=1.662
cc_201 VPB N_A_1034_368#_c_843_n 0.0172781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1367_92#_c_1044_n 0.0227981f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_203 VPB N_A_1367_92#_c_1045_n 0.0211965f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_204 VPB N_A_1367_92#_c_1038_n 0.00197089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_1367_92#_c_1039_n 0.0231488f $X=-0.19 $Y=1.66 $X2=2.395 $Y2=1.575
cc_206 VPB N_A_1367_92#_c_1048_n 0.00178601f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.575
cc_207 VPB N_A_1367_92#_c_1049_n 0.00224162f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_208 VPB N_A_1367_92#_c_1043_n 0.00122099f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.67
cc_209 VPB N_A_1233_118#_c_1147_n 0.0164911f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_210 VPB N_A_1233_118#_c_1156_n 0.015497f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_211 VPB N_A_1233_118#_c_1157_n 5.61498e-19 $X=-0.19 $Y=1.66 $X2=2.395
+ $Y2=1.575
cc_212 VPB N_A_1233_118#_c_1149_n 0.00734892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1233_118#_c_1150_n 0.0125171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1233_118#_c_1153_n 0.00754174f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.67
cc_215 VPB N_A_1233_118#_c_1161_n 0.00112616f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.26
cc_216 VPB N_A_855_368#_c_1280_n 0.0226181f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_217 VPB N_A_855_368#_c_1283_n 0.0774298f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_218 VPB N_A_855_368#_c_1298_n 0.0597393f $X=-0.19 $Y=1.66 $X2=2.395 $Y2=1.575
cc_219 VPB N_A_855_368#_c_1299_n 0.0123764f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.575
cc_220 VPB N_A_855_368#_c_1300_n 0.00781624f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.575
cc_221 VPB N_A_855_368#_c_1301_n 0.0174462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_855_368#_c_1302_n 0.0159175f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_223 VPB N_A_855_368#_c_1303_n 0.187923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_855_368#_c_1304_n 0.0078517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_855_368#_c_1305_n 0.0132688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_855_368#_M1004_g 0.00887153f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_227 VPB N_A_855_368#_c_1286_n 0.0193138f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_228 VPB N_A_855_368#_c_1287_n 0.00438317f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_229 VPB N_A_855_368#_c_1309_n 0.0089865f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.662
cc_230 VPB N_A_855_368#_c_1310_n 0.00271787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_855_368#_c_1294_n 0.00279634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_855_368#_c_1312_n 0.00185216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1997_272#_c_1483_n 0.0211446f $X=-0.19 $Y=1.66 $X2=1.005
+ $Y2=2.155
cc_234 VPB N_A_1997_272#_c_1494_n 0.0298064f $X=-0.19 $Y=1.66 $X2=1.005
+ $Y2=2.245
cc_235 VPB N_A_1997_272#_c_1495_n 0.0223998f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_236 VPB N_A_1997_272#_c_1496_n 0.00909249f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_237 VPB N_A_1997_272#_c_1491_n 0.00705302f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_238 VPB N_A_1745_74#_c_1600_n 0.00901615f $X=-0.19 $Y=1.66 $X2=1.005
+ $Y2=2.245
cc_239 VPB N_A_1745_74#_c_1611_n 0.0207522f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_240 VPB N_A_1745_74#_c_1612_n 0.0222832f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=1.26
cc_241 VPB N_A_1745_74#_c_1613_n 0.0425889f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.575
cc_242 VPB N_A_1745_74#_c_1614_n 0.018388f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.425
cc_243 VPB N_A_1745_74#_c_1615_n 0.00552913f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_244 VPB N_A_1745_74#_c_1616_n 0.00178486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1745_74#_c_1605_n 0.00223832f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_246 VPB N_A_1745_74#_c_1618_n 0.00730775f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.425
cc_247 VPB N_A_1745_74#_c_1619_n 0.00277122f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.26
cc_248 VPB N_A_1745_74#_c_1620_n 0.00536408f $X=-0.19 $Y=1.66 $X2=1.623
+ $Y2=1.662
cc_249 VPB N_A_2399_424#_c_1771_n 0.021165f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_250 VPB N_A_2399_424#_c_1767_n 0.00855036f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=1.26
cc_251 VPB N_A_2399_424#_c_1773_n 0.0138904f $X=-0.19 $Y=1.66 $X2=2.395
+ $Y2=1.575
cc_252 VPB N_A_2399_424#_c_1769_n 0.0133083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1814_n 0.00651803f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_254 VPB N_VPWR_c_1815_n 0.00662228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1816_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.67
cc_256 VPB N_VPWR_c_1817_n 0.0144445f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_257 VPB N_VPWR_c_1818_n 0.02311f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.26
cc_258 VPB N_VPWR_c_1819_n 0.0144685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1820_n 0.0127921f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.662
cc_260 VPB N_VPWR_c_1821_n 0.0158276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1822_n 0.0193772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1823_n 0.0379482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1824_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1825_n 0.0523435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1826_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1827_n 0.020808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1828_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1829_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1830_n 0.0596953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1831_n 0.0636234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1832_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1833_n 0.0181474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1813_n 0.127682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1835_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1836_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1837_n 0.00443527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1838_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1839_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_300_464#_c_1982_n 0.00671604f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_280 VPB N_A_300_464#_c_1976_n 0.00482108f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.575
cc_281 VPB N_A_300_464#_c_1984_n 0.0125755f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_282 VPB N_A_300_464#_c_1985_n 0.00122623f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_283 VPB N_A_300_464#_c_1986_n 0.00285414f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.67
cc_284 VPB N_A_300_464#_c_1987_n 0.00709116f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_285 VPB N_A_300_464#_c_1988_n 0.00193082f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_286 VPB N_A_300_464#_c_1980_n 0.00530725f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.26
cc_287 VPB N_A_300_464#_c_1990_n 0.00267737f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.662
cc_288 VPB N_A_300_464#_c_1991_n 0.00929993f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.665
cc_289 VPB Q 0.0544732f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_290 N_SCE_M1037_g N_A_27_88#_c_379_n 0.00834942f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_291 N_SCE_M1037_g N_A_27_88#_c_380_n 0.0131974f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_292 N_SCE_c_296_n N_A_27_88#_c_380_n 0.0103131f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_293 N_SCE_c_297_n N_A_27_88#_c_380_n 0.0273678f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_294 N_SCE_c_299_n N_A_27_88#_c_387_n 0.0130468f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_295 N_SCE_c_301_n N_A_27_88#_c_387_n 8.82207e-19 $X=1.005 $Y=2.245 $X2=0
+ $Y2=0
cc_296 N_SCE_M1037_g N_A_27_88#_c_381_n 0.0204376f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_297 N_SCE_c_296_n N_A_27_88#_c_381_n 0.0032453f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_298 N_SCE_c_297_n N_A_27_88#_c_381_n 0.0382971f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_299 N_SCE_c_293_n N_A_27_88#_c_388_n 0.0271109f $X=2.395 $Y=1.575 $X2=0 $Y2=0
cc_300 N_SCE_c_294_n N_A_27_88#_c_389_n 0.0249956f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_301 N_SCE_c_295_n N_A_27_88#_c_389_n 3.39021e-19 $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_302 N_SCE_c_293_n N_A_27_88#_c_390_n 0.00722834f $X=2.395 $Y=1.575 $X2=0
+ $Y2=0
cc_303 N_SCE_c_294_n N_A_27_88#_c_390_n 0.00200458f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_304 N_SCE_c_295_n N_A_27_88#_c_390_n 0.016847f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_305 N_SCE_c_298_n N_A_27_88#_c_391_n 0.00495347f $X=0.505 $Y=2.155 $X2=0
+ $Y2=0
cc_306 N_SCE_c_299_n N_A_27_88#_c_391_n 4.59028e-19 $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_307 N_SCE_M1037_g N_A_27_88#_c_383_n 7.61834e-19 $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_308 N_SCE_c_297_n N_A_27_88#_c_383_n 0.0212113f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_309 N_SCE_M1037_g N_A_27_88#_c_384_n 0.00727818f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_310 N_SCE_c_296_n N_A_27_88#_c_384_n 0.00441678f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_311 N_SCE_c_297_n N_A_27_88#_c_384_n 0.008287f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_312 N_SCE_c_298_n N_A_27_88#_c_392_n 0.00636452f $X=0.505 $Y=2.155 $X2=0
+ $Y2=0
cc_313 N_SCE_c_299_n N_A_27_88#_c_392_n 0.00700767f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_314 N_SCE_c_300_n N_A_27_88#_c_392_n 0.00899514f $X=1.005 $Y=2.155 $X2=0
+ $Y2=0
cc_315 N_SCE_c_301_n N_A_27_88#_c_392_n 0.007641f $X=1.005 $Y=2.245 $X2=0 $Y2=0
cc_316 N_SCE_c_293_n N_A_27_88#_c_392_n 0.0110297f $X=2.395 $Y=1.575 $X2=0 $Y2=0
cc_317 N_SCE_c_296_n N_A_27_88#_c_392_n 0.00381149f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_318 N_SCE_c_297_n N_A_27_88#_c_392_n 0.101415f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_319 N_SCE_c_301_n N_D_c_468_n 0.0373647f $X=1.005 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_320 N_SCE_c_300_n N_D_c_462_n 0.0062192f $X=1.005 $Y=2.155 $X2=0 $Y2=0
cc_321 N_SCE_c_297_n N_D_c_462_n 0.00447951f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_322 N_SCE_c_305_n N_D_c_462_n 0.00931586f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_323 N_SCE_c_294_n N_D_c_463_n 0.00125287f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_324 N_SCE_c_295_n N_D_c_463_n 0.00839725f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_325 N_SCE_c_300_n N_D_c_470_n 0.0098871f $X=1.005 $Y=2.155 $X2=0 $Y2=0
cc_326 N_SCE_c_297_n N_D_c_470_n 0.00173212f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_327 N_SCE_c_293_n N_D_c_464_n 0.00669247f $X=2.395 $Y=1.575 $X2=0 $Y2=0
cc_328 N_SCE_c_296_n N_D_c_464_n 0.00663484f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_329 N_SCE_c_297_n N_D_c_464_n 0.00195725f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_330 N_SCE_c_305_n N_D_c_464_n 0.0037388f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_331 N_SCE_M1030_g N_D_c_465_n 0.00676226f $X=2.65 $Y=0.615 $X2=0 $Y2=0
cc_332 N_SCE_c_293_n N_D_c_465_n 0.00318874f $X=2.395 $Y=1.575 $X2=0 $Y2=0
cc_333 N_SCE_c_295_n N_D_c_465_n 2.48719e-19 $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_334 N_SCE_M1030_g N_D_c_466_n 0.00133517f $X=2.65 $Y=0.615 $X2=0 $Y2=0
cc_335 N_SCE_c_297_n N_D_c_466_n 0.0338107f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_336 N_SCE_M1030_g N_D_c_467_n 0.00735939f $X=2.65 $Y=0.615 $X2=0 $Y2=0
cc_337 N_SCE_M1030_g N_SCD_M1021_g 0.0632491f $X=2.65 $Y=0.615 $X2=0 $Y2=0
cc_338 N_SCE_c_294_n N_SCD_M1021_g 0.00116379f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_339 N_SCE_c_294_n SCD 0.0136985f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_340 N_SCE_c_295_n SCD 5.33056e-19 $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_341 N_SCE_c_294_n N_SCD_c_519_n 0.00206106f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_342 N_SCE_c_295_n N_SCD_c_519_n 0.00863742f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_343 N_SCE_c_299_n N_VPWR_c_1814_n 0.00657693f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_344 N_SCE_c_301_n N_VPWR_c_1814_n 0.0146782f $X=1.005 $Y=2.245 $X2=0 $Y2=0
cc_345 N_SCE_c_299_n N_VPWR_c_1829_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_346 N_SCE_c_301_n N_VPWR_c_1830_n 0.00413917f $X=1.005 $Y=2.245 $X2=0 $Y2=0
cc_347 N_SCE_c_299_n N_VPWR_c_1813_n 0.00860873f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_348 N_SCE_c_301_n N_VPWR_c_1813_n 0.00817532f $X=1.005 $Y=2.245 $X2=0 $Y2=0
cc_349 N_SCE_c_301_n N_A_300_464#_c_1982_n 0.00181955f $X=1.005 $Y=2.245 $X2=0
+ $Y2=0
cc_350 N_SCE_M1030_g N_A_300_464#_c_1975_n 0.00897301f $X=2.65 $Y=0.615 $X2=0
+ $Y2=0
cc_351 N_SCE_c_294_n N_A_300_464#_c_1975_n 0.00904054f $X=2.56 $Y=1.425 $X2=0
+ $Y2=0
cc_352 N_SCE_M1030_g N_A_300_464#_c_1981_n 0.0111649f $X=2.65 $Y=0.615 $X2=0
+ $Y2=0
cc_353 N_SCE_c_293_n N_A_300_464#_c_1981_n 0.00563615f $X=2.395 $Y=1.575 $X2=0
+ $Y2=0
cc_354 N_SCE_c_294_n N_A_300_464#_c_1981_n 0.016885f $X=2.56 $Y=1.425 $X2=0
+ $Y2=0
cc_355 N_SCE_c_295_n N_A_300_464#_c_1981_n 0.0013723f $X=2.56 $Y=1.425 $X2=0
+ $Y2=0
cc_356 N_SCE_M1037_g N_VGND_c_2147_n 0.0142996f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_357 N_SCE_M1030_g N_VGND_c_2153_n 9.15902e-19 $X=2.65 $Y=0.615 $X2=0 $Y2=0
cc_358 N_SCE_M1037_g N_VGND_c_2157_n 0.00438299f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_359 N_SCE_M1037_g N_VGND_c_2163_n 0.00439883f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_360 N_SCE_M1030_g N_noxref_24_c_2273_n 0.0133411f $X=2.65 $Y=0.615 $X2=0
+ $Y2=0
cc_361 N_SCE_M1037_g N_noxref_24_c_2274_n 8.90151e-19 $X=0.495 $Y=0.65 $X2=0
+ $Y2=0
cc_362 N_A_27_88#_c_388_n N_D_c_462_n 0.0010716f $X=2.207 $Y=2.002 $X2=0 $Y2=0
cc_363 N_A_27_88#_c_390_n N_D_c_462_n 0.0150513f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_364 N_A_27_88#_c_392_n N_D_c_462_n 0.00500376f $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_365 N_A_27_88#_c_392_n N_D_c_470_n 0.0191365f $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_366 N_A_27_88#_c_392_n N_D_c_464_n 7.9327e-19 $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_367 N_A_27_88#_c_390_n N_D_c_465_n 9.15182e-19 $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_368 N_A_27_88#_c_383_n N_D_c_465_n 2.69613e-19 $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_369 N_A_27_88#_c_384_n N_D_c_465_n 0.0143534f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_370 N_A_27_88#_c_378_n N_D_c_466_n 0.00484268f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_371 N_A_27_88#_c_383_n N_D_c_466_n 0.0250153f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_372 N_A_27_88#_c_384_n N_D_c_466_n 0.0014755f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_373 N_A_27_88#_c_378_n N_D_c_467_n 0.0356736f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_374 N_A_27_88#_c_385_n N_SCD_c_520_n 0.0390364f $X=2.615 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_375 N_A_27_88#_c_385_n N_SCD_c_517_n 0.0225329f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_376 N_A_27_88#_c_389_n N_SCD_c_517_n 0.00131024f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_377 N_A_27_88#_c_385_n SCD 4.03756e-19 $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_378 N_A_27_88#_c_389_n SCD 0.019263f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_379 N_A_27_88#_c_387_n N_VPWR_c_1814_n 0.0246172f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_380 N_A_27_88#_c_392_n N_VPWR_c_1814_n 0.0234317f $X=2.035 $Y=2.002 $X2=0
+ $Y2=0
cc_381 N_A_27_88#_c_385_n N_VPWR_c_1815_n 0.00139568f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_382 N_A_27_88#_c_387_n N_VPWR_c_1829_n 0.0145938f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_383 N_A_27_88#_c_385_n N_VPWR_c_1830_n 0.00444483f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_384 N_A_27_88#_c_385_n N_VPWR_c_1813_n 0.0045343f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_385 N_A_27_88#_c_387_n N_VPWR_c_1813_n 0.0120466f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_386 N_A_27_88#_c_390_n N_A_300_464#_c_1982_n 0.00356798f $X=2.54 $Y=1.995
+ $X2=0 $Y2=0
cc_387 N_A_27_88#_c_392_n N_A_300_464#_c_1982_n 0.0311708f $X=2.035 $Y=2.002
+ $X2=0 $Y2=0
cc_388 N_A_27_88#_c_385_n N_A_300_464#_c_2001_n 0.00887275f $X=2.615 $Y=2.245
+ $X2=0 $Y2=0
cc_389 N_A_27_88#_c_389_n N_A_300_464#_c_2001_n 0.0311708f $X=2.54 $Y=1.995
+ $X2=0 $Y2=0
cc_390 N_A_27_88#_c_385_n N_A_300_464#_c_1990_n 0.00919805f $X=2.615 $Y=2.245
+ $X2=0 $Y2=0
cc_391 N_A_27_88#_c_388_n N_A_300_464#_c_1990_n 0.0311708f $X=2.207 $Y=2.002
+ $X2=0 $Y2=0
cc_392 N_A_27_88#_c_378_n N_VGND_c_2147_n 0.00578639f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_393 N_A_27_88#_c_379_n N_VGND_c_2147_n 0.0179429f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_394 N_A_27_88#_c_381_n N_VGND_c_2147_n 0.0279517f $X=1.045 $Y=1.157 $X2=0
+ $Y2=0
cc_395 N_A_27_88#_c_378_n N_VGND_c_2153_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_396 N_A_27_88#_c_379_n N_VGND_c_2157_n 0.00862619f $X=0.28 $Y=0.65 $X2=0
+ $Y2=0
cc_397 N_A_27_88#_c_379_n N_VGND_c_2163_n 0.00876292f $X=0.28 $Y=0.65 $X2=0
+ $Y2=0
cc_398 N_A_27_88#_c_378_n N_noxref_24_c_2273_n 0.0108727f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_399 N_A_27_88#_c_378_n N_noxref_24_c_2274_n 0.00859442f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_400 N_A_27_88#_c_383_n N_noxref_24_c_2274_n 0.0133426f $X=1.21 $Y=1.1 $X2=0
+ $Y2=0
cc_401 N_A_27_88#_c_384_n N_noxref_24_c_2274_n 0.0017694f $X=1.21 $Y=1.1 $X2=0
+ $Y2=0
cc_402 N_D_c_468_n N_VPWR_c_1814_n 0.00237824f $X=1.425 $Y=2.245 $X2=0 $Y2=0
cc_403 N_D_c_468_n N_VPWR_c_1830_n 0.00444483f $X=1.425 $Y=2.245 $X2=0 $Y2=0
cc_404 N_D_c_468_n N_VPWR_c_1813_n 0.00859301f $X=1.425 $Y=2.245 $X2=0 $Y2=0
cc_405 N_D_c_466_n N_A_300_464#_M1013_d 0.00160189f $X=1.935 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_406 N_D_c_468_n N_A_300_464#_c_1982_n 0.0115052f $X=1.425 $Y=2.245 $X2=0
+ $Y2=0
cc_407 N_D_c_470_n N_A_300_464#_c_1982_n 0.00629416f $X=1.425 $Y=2.16 $X2=0
+ $Y2=0
cc_408 N_D_c_465_n N_A_300_464#_c_1981_n 6.29158e-19 $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_409 N_D_c_466_n N_A_300_464#_c_1981_n 0.0234916f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_410 N_D_c_467_n N_A_300_464#_c_1981_n 0.00518029f $X=1.935 $Y=0.935 $X2=0
+ $Y2=0
cc_411 N_D_c_467_n N_VGND_c_2153_n 9.15902e-19 $X=1.935 $Y=0.935 $X2=0 $Y2=0
cc_412 N_D_c_465_n N_noxref_24_c_2273_n 5.66605e-19 $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_413 N_D_c_466_n N_noxref_24_c_2273_n 0.0128576f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_414 N_D_c_467_n N_noxref_24_c_2273_n 0.011902f $X=1.935 $Y=0.935 $X2=0 $Y2=0
cc_415 N_D_c_467_n N_noxref_24_c_2274_n 0.00113655f $X=1.935 $Y=0.935 $X2=0
+ $Y2=0
cc_416 N_D_c_466_n noxref_25 0.00198619f $X=1.935 $Y=1.1 $X2=-0.19 $Y2=-0.245
cc_417 N_SCD_c_520_n N_RESET_B_c_568_n 0.0163314f $X=3.035 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_418 N_SCD_c_517_n N_RESET_B_c_568_n 0.0198798f $X=3.11 $Y=1.945 $X2=-0.19
+ $Y2=-0.245
cc_419 SCD N_RESET_B_c_568_n 2.37625e-19 $X=3.035 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_420 N_SCD_M1021_g N_RESET_B_M1016_g 0.0267916f $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_421 SCD N_RESET_B_M1016_g 5.82635e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_422 N_SCD_c_519_n N_RESET_B_M1016_g 0.0108821f $X=3.11 $Y=1.605 $X2=0 $Y2=0
cc_423 N_SCD_c_520_n N_VPWR_c_1815_n 0.00912975f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_424 N_SCD_c_520_n N_VPWR_c_1830_n 0.00413917f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_425 N_SCD_c_520_n N_VPWR_c_1813_n 0.00408655f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_426 N_SCD_c_520_n N_A_300_464#_c_2001_n 0.0123812f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_427 N_SCD_c_517_n N_A_300_464#_c_2001_n 8.1818e-19 $X=3.11 $Y=1.945 $X2=0
+ $Y2=0
cc_428 SCD N_A_300_464#_c_2001_n 0.0212424f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_429 N_SCD_M1021_g N_A_300_464#_c_1975_n 0.013373f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_430 SCD N_A_300_464#_c_1975_n 0.0146824f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_431 N_SCD_c_519_n N_A_300_464#_c_1975_n 0.00106413f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_432 N_SCD_c_520_n N_A_300_464#_c_1976_n 0.00151656f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_433 N_SCD_M1021_g N_A_300_464#_c_1976_n 0.00645124f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_434 N_SCD_c_517_n N_A_300_464#_c_1976_n 0.00183512f $X=3.11 $Y=1.945 $X2=0
+ $Y2=0
cc_435 SCD N_A_300_464#_c_1976_n 0.0534507f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_436 N_SCD_c_519_n N_A_300_464#_c_1976_n 0.00426807f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_437 N_SCD_c_520_n N_A_300_464#_c_1985_n 5.39484e-19 $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_438 N_SCD_c_520_n N_A_300_464#_c_1990_n 0.00165456f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_439 N_SCD_M1021_g N_A_300_464#_c_1981_n 0.00143504f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_440 N_SCD_c_520_n N_A_300_464#_c_1991_n 4.29898e-19 $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_441 N_SCD_M1021_g N_VGND_c_2153_n 9.09582e-19 $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_442 N_SCD_M1021_g N_noxref_24_c_2273_n 0.0226823f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_443 N_RESET_B_c_575_n N_CLK_c_772_n 0.00217906f $X=7.775 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_444 N_RESET_B_c_581_n N_CLK_c_772_n 0.0039069f $X=3.95 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_445 N_RESET_B_c_582_n N_CLK_c_772_n 4.10166e-19 $X=3.95 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_446 N_RESET_B_M1016_g N_CLK_c_774_n 0.016727f $X=3.655 $Y=0.615 $X2=0 $Y2=0
cc_447 N_RESET_B_c_575_n N_CLK_c_774_n 0.00236558f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_448 N_RESET_B_c_576_n N_CLK_c_774_n 0.00141283f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_449 N_RESET_B_c_581_n N_CLK_c_774_n 0.00750615f $X=3.95 $Y=1.995 $X2=0 $Y2=0
cc_450 N_RESET_B_c_582_n N_CLK_c_774_n 0.00162476f $X=3.95 $Y=1.995 $X2=0 $Y2=0
cc_451 N_RESET_B_c_575_n N_CLK_c_785_n 0.0055905f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_452 N_RESET_B_M1016_g N_CLK_c_775_n 0.00407861f $X=3.655 $Y=0.615 $X2=0 $Y2=0
cc_453 N_RESET_B_c_576_n N_CLK_c_775_n 0.00358597f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_454 N_RESET_B_c_581_n N_CLK_c_775_n 6.43181e-19 $X=3.95 $Y=1.995 $X2=0 $Y2=0
cc_455 N_RESET_B_c_582_n N_CLK_c_775_n 0.0104674f $X=3.95 $Y=1.995 $X2=0 $Y2=0
cc_456 N_RESET_B_c_575_n N_A_1034_368#_c_845_n 0.00340123f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_457 N_RESET_B_c_575_n N_A_1034_368#_c_824_n 0.0039938f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_458 N_RESET_B_c_577_n N_A_1034_368#_c_848_n 0.00642678f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_459 N_RESET_B_c_575_n N_A_1034_368#_c_832_n 0.0355245f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_460 N_RESET_B_c_575_n N_A_1034_368#_c_833_n 0.0164707f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_461 N_RESET_B_c_561_n N_A_1034_368#_c_834_n 0.0029615f $X=7.3 $Y=1.085 $X2=0
+ $Y2=0
cc_462 N_RESET_B_c_561_n N_A_1034_368#_c_835_n 0.0119788f $X=7.3 $Y=1.085 $X2=0
+ $Y2=0
cc_463 N_RESET_B_c_562_n N_A_1034_368#_c_835_n 0.0016592f $X=7.595 $Y=1.16 $X2=0
+ $Y2=0
cc_464 N_RESET_B_c_561_n N_A_1034_368#_c_862_n 0.00273826f $X=7.3 $Y=1.085 $X2=0
+ $Y2=0
cc_465 N_RESET_B_c_577_n N_A_1034_368#_c_839_n 0.0173785f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_466 N_RESET_B_c_577_n N_A_1034_368#_c_852_n 0.0197423f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_467 N_RESET_B_c_575_n N_A_1034_368#_c_843_n 0.00379596f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_468 N_RESET_B_c_577_n N_A_1367_92#_M1001_d 0.00464147f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_469 N_RESET_B_c_561_n N_A_1367_92#_M1027_g 0.0386216f $X=7.3 $Y=1.085 $X2=0
+ $Y2=0
cc_470 N_RESET_B_c_564_n N_A_1367_92#_M1027_g 0.00277736f $X=7.67 $Y=1.815 $X2=0
+ $Y2=0
cc_471 N_RESET_B_c_564_n N_A_1367_92#_c_1044_n 0.00501376f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_472 N_RESET_B_c_575_n N_A_1367_92#_c_1044_n 0.0101236f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_473 N_RESET_B_c_571_n N_A_1367_92#_c_1045_n 0.01292f $X=7.685 $Y=2.23 $X2=0
+ $Y2=0
cc_474 N_RESET_B_c_583_n N_A_1367_92#_c_1045_n 0.00501376f $X=7.685 $Y=2.022
+ $X2=0 $Y2=0
cc_475 N_RESET_B_c_563_n N_A_1367_92#_c_1038_n 0.00963889f $X=7.375 $Y=1.16
+ $X2=0 $Y2=0
cc_476 N_RESET_B_c_564_n N_A_1367_92#_c_1038_n 0.00161804f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_477 N_RESET_B_c_575_n N_A_1367_92#_c_1038_n 0.00823427f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_478 N_RESET_B_c_563_n N_A_1367_92#_c_1039_n 0.00715091f $X=7.375 $Y=1.16
+ $X2=0 $Y2=0
cc_479 N_RESET_B_c_564_n N_A_1367_92#_c_1039_n 0.0173421f $X=7.67 $Y=1.815 $X2=0
+ $Y2=0
cc_480 N_RESET_B_c_575_n N_A_1367_92#_c_1039_n 0.00318126f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_481 N_RESET_B_c_561_n N_A_1367_92#_c_1040_n 0.00534949f $X=7.3 $Y=1.085 $X2=0
+ $Y2=0
cc_482 N_RESET_B_c_562_n N_A_1367_92#_c_1040_n 0.0141377f $X=7.595 $Y=1.16 $X2=0
+ $Y2=0
cc_483 N_RESET_B_c_563_n N_A_1367_92#_c_1040_n 0.00131223f $X=7.375 $Y=1.16
+ $X2=0 $Y2=0
cc_484 N_RESET_B_c_561_n N_A_1367_92#_c_1041_n 0.00414754f $X=7.3 $Y=1.085 $X2=0
+ $Y2=0
cc_485 N_RESET_B_c_577_n N_A_1367_92#_c_1049_n 0.0360053f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_486 N_RESET_B_c_562_n N_A_1233_118#_M1033_g 0.00636759f $X=7.595 $Y=1.16
+ $X2=0 $Y2=0
cc_487 N_RESET_B_c_577_n N_A_1233_118#_c_1147_n 3.01246e-19 $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_488 N_RESET_B_c_577_n N_A_1233_118#_c_1156_n 0.0082395f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_489 N_RESET_B_c_575_n N_A_1233_118#_c_1157_n 0.00861368f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_490 N_RESET_B_c_561_n N_A_1233_118#_c_1148_n 3.96747e-19 $X=7.3 $Y=1.085
+ $X2=0 $Y2=0
cc_491 N_RESET_B_c_575_n N_A_1233_118#_c_1149_n 0.0240634f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_492 N_RESET_B_c_575_n N_A_1233_118#_c_1168_n 0.0215639f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_493 N_RESET_B_c_564_n N_A_1233_118#_c_1150_n 0.0113497f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_494 N_RESET_B_c_571_n N_A_1233_118#_c_1150_n 0.0182508f $X=7.685 $Y=2.23
+ $X2=0 $Y2=0
cc_495 N_RESET_B_c_575_n N_A_1233_118#_c_1150_n 0.0273088f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_496 N_RESET_B_c_578_n N_A_1233_118#_c_1150_n 0.01197f $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_497 N_RESET_B_c_579_n N_A_1233_118#_c_1150_n 0.0389238f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_498 N_RESET_B_c_583_n N_A_1233_118#_c_1150_n 0.0165391f $X=7.685 $Y=2.022
+ $X2=0 $Y2=0
cc_499 N_RESET_B_c_562_n N_A_1233_118#_c_1151_n 0.0023739f $X=7.595 $Y=1.16
+ $X2=0 $Y2=0
cc_500 N_RESET_B_c_564_n N_A_1233_118#_c_1151_n 0.00614229f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_501 N_RESET_B_c_564_n N_A_1233_118#_c_1152_n 0.00830382f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_502 N_RESET_B_c_575_n N_A_1233_118#_c_1152_n 0.00357593f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_503 N_RESET_B_c_577_n N_A_1233_118#_c_1152_n 0.00581394f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_504 N_RESET_B_c_578_n N_A_1233_118#_c_1152_n 0.00371961f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_505 N_RESET_B_c_579_n N_A_1233_118#_c_1152_n 0.0172409f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_506 N_RESET_B_c_583_n N_A_1233_118#_c_1152_n 0.00735754f $X=7.685 $Y=2.022
+ $X2=0 $Y2=0
cc_507 N_RESET_B_c_564_n N_A_1233_118#_c_1153_n 0.0188449f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_508 N_RESET_B_c_577_n N_A_1233_118#_c_1153_n 0.00593186f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_509 N_RESET_B_c_579_n N_A_1233_118#_c_1153_n 6.74459e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_510 N_RESET_B_c_583_n N_A_1233_118#_c_1153_n 0.0093828f $X=7.685 $Y=2.022
+ $X2=0 $Y2=0
cc_511 N_RESET_B_c_575_n N_A_855_368#_M1022_s 0.0011702f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_512 N_RESET_B_c_575_n N_A_855_368#_c_1280_n 0.00478768f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_513 N_RESET_B_c_575_n N_A_855_368#_c_1283_n 0.0023679f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_514 N_RESET_B_c_575_n N_A_855_368#_c_1302_n 0.00394165f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_515 N_RESET_B_c_571_n N_A_855_368#_c_1303_n 0.00949691f $X=7.685 $Y=2.23
+ $X2=0 $Y2=0
cc_516 N_RESET_B_c_577_n N_A_855_368#_M1004_g 0.0137675f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_517 N_RESET_B_c_577_n N_A_855_368#_c_1286_n 0.00383889f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_518 N_RESET_B_c_577_n N_A_855_368#_c_1287_n 2.83807e-19 $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_519 N_RESET_B_M1016_g N_A_855_368#_c_1292_n 0.00433927f $X=3.655 $Y=0.615
+ $X2=0 $Y2=0
cc_520 N_RESET_B_M1016_g N_A_855_368#_c_1322_n 0.00423005f $X=3.655 $Y=0.615
+ $X2=0 $Y2=0
cc_521 N_RESET_B_c_575_n N_A_855_368#_c_1310_n 0.0156654f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_522 N_RESET_B_c_568_n N_A_855_368#_c_1312_n 0.00134964f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_523 N_RESET_B_M1016_g N_A_855_368#_c_1312_n 2.17516e-19 $X=3.655 $Y=0.615
+ $X2=0 $Y2=0
cc_524 N_RESET_B_c_575_n N_A_855_368#_c_1312_n 0.014404f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_525 N_RESET_B_c_576_n N_A_855_368#_c_1312_n 0.00277564f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_526 N_RESET_B_c_581_n N_A_855_368#_c_1312_n 0.00101677f $X=3.95 $Y=1.995
+ $X2=0 $Y2=0
cc_527 N_RESET_B_c_582_n N_A_855_368#_c_1312_n 0.0240037f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_528 N_RESET_B_c_575_n N_A_855_368#_c_1295_n 0.00730094f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_529 N_RESET_B_M1038_g N_A_1997_272#_M1005_g 0.0312551f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_530 N_RESET_B_c_566_n N_A_1997_272#_c_1483_n 0.0225363f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_531 N_RESET_B_c_567_n N_A_1997_272#_c_1483_n 0.00643996f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_532 N_RESET_B_c_584_n N_A_1997_272#_c_1483_n 0.00119422f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_573_n N_A_1997_272#_c_1494_n 0.00511887f $X=10.885 $Y=2.375
+ $X2=0 $Y2=0
cc_534 N_RESET_B_c_577_n N_A_1997_272#_c_1494_n 0.00508273f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_535 N_RESET_B_c_585_n N_A_1997_272#_c_1494_n 0.0128577f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_536 N_RESET_B_c_574_n N_A_1997_272#_c_1495_n 0.0138023f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_537 N_RESET_B_c_566_n N_A_1997_272#_c_1484_n 0.00935059f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_567_n N_A_1997_272#_c_1484_n 0.0053082f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_539 RESET_B N_A_1997_272#_c_1484_n 0.00164136f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_540 N_RESET_B_c_584_n N_A_1997_272#_c_1484_n 0.0191591f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_541 N_RESET_B_c_585_n N_A_1997_272#_c_1484_n 0.00143438f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_542 N_RESET_B_M1038_g N_A_1997_272#_c_1485_n 0.00111706f $X=10.6 $Y=0.58
+ $X2=0 $Y2=0
cc_543 N_RESET_B_M1038_g N_A_1997_272#_c_1488_n 7.22053e-19 $X=10.6 $Y=0.58
+ $X2=0 $Y2=0
cc_544 N_RESET_B_c_577_n N_A_1997_272#_c_1490_n 0.0131744f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_574_n N_A_1997_272#_c_1496_n 0.00680136f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_584_n N_A_1997_272#_c_1496_n 9.92047e-19 $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_566_n N_A_1997_272#_c_1491_n 0.00366777f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_574_n N_A_1997_272#_c_1491_n 0.00111437f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_549 RESET_B N_A_1997_272#_c_1491_n 0.00158814f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_550 N_RESET_B_c_584_n N_A_1997_272#_c_1491_n 0.0232461f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_551 N_RESET_B_c_585_n N_A_1997_272#_c_1491_n 0.00858202f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_552 N_RESET_B_c_577_n N_A_1745_74#_M1004_d 0.00297016f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_553 N_RESET_B_M1038_g N_A_1745_74#_M1028_g 0.0518692f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_567_n N_A_1745_74#_c_1600_n 0.0117915f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_584_n N_A_1745_74#_c_1600_n 3.43698e-19 $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_556 N_RESET_B_c_585_n N_A_1745_74#_c_1600_n 0.00946465f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_557 N_RESET_B_c_574_n N_A_1745_74#_c_1611_n 0.00946465f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_558 N_RESET_B_c_574_n N_A_1745_74#_c_1612_n 0.00921795f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_559 N_RESET_B_M1038_g N_A_1745_74#_c_1602_n 0.00646231f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_567_n N_A_1745_74#_c_1602_n 0.0030434f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_573_n N_A_1745_74#_c_1615_n 0.00946465f $X=10.885 $Y=2.375
+ $X2=0 $Y2=0
cc_562 N_RESET_B_c_577_n N_A_1745_74#_c_1616_n 0.00561127f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_563 N_RESET_B_c_566_n N_A_1745_74#_c_1618_n 6.20198e-19 $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_564 N_RESET_B_c_577_n N_A_1745_74#_c_1618_n 0.0131083f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_565 RESET_B N_A_1745_74#_c_1618_n 2.51275e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_566 N_RESET_B_c_584_n N_A_1745_74#_c_1618_n 0.00608543f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_567 N_RESET_B_c_577_n N_A_1745_74#_c_1619_n 0.0053742f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_568 N_RESET_B_c_573_n N_A_1745_74#_c_1620_n 0.00159843f $X=10.885 $Y=2.375
+ $X2=0 $Y2=0
cc_569 N_RESET_B_c_574_n N_A_1745_74#_c_1620_n 2.78257e-19 $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_570 N_RESET_B_c_577_n N_A_1745_74#_c_1620_n 0.020931f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_571 RESET_B N_A_1745_74#_c_1620_n 3.29892e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_572 N_RESET_B_c_584_n N_A_1745_74#_c_1620_n 0.00622512f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_573 N_RESET_B_c_585_n N_A_1745_74#_c_1620_n 6.08738e-19 $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_574 N_RESET_B_M1038_g N_A_1745_74#_c_1609_n 0.015752f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_567_n N_A_1745_74#_c_1609_n 0.00357206f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_576 N_RESET_B_c_575_n N_VPWR_M1022_d 0.0030901f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_577 N_RESET_B_c_577_n N_VPWR_M1001_s 0.00689173f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_568_n N_VPWR_c_1815_n 0.00571347f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_579 N_RESET_B_c_571_n N_VPWR_c_1817_n 0.00404752f $X=7.685 $Y=2.23 $X2=0
+ $Y2=0
cc_580 N_RESET_B_c_575_n N_VPWR_c_1817_n 7.58628e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_581 N_RESET_B_c_564_n N_VPWR_c_1819_n 0.00146391f $X=7.67 $Y=1.815 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_571_n N_VPWR_c_1819_n 0.00504716f $X=7.685 $Y=2.23 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_577_n N_VPWR_c_1819_n 0.0185404f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_584 N_RESET_B_c_578_n N_VPWR_c_1819_n 5.19261e-19 $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_585 N_RESET_B_c_579_n N_VPWR_c_1819_n 0.0183634f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_586 N_RESET_B_c_583_n N_VPWR_c_1819_n 0.00295171f $X=7.685 $Y=2.022 $X2=0
+ $Y2=0
cc_587 N_RESET_B_c_574_n N_VPWR_c_1820_n 0.00720194f $X=10.885 $Y=2.465 $X2=0
+ $Y2=0
cc_588 N_RESET_B_c_577_n N_VPWR_c_1820_n 0.00652534f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_589 RESET_B N_VPWR_c_1820_n 6.45709e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_590 N_RESET_B_c_584_n N_VPWR_c_1820_n 0.00292772f $X=10.805 $Y=1.985 $X2=0
+ $Y2=0
cc_591 N_RESET_B_c_585_n N_VPWR_c_1820_n 6.5955e-19 $X=10.885 $Y=1.985 $X2=0
+ $Y2=0
cc_592 N_RESET_B_c_568_n N_VPWR_c_1823_n 0.00445602f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_574_n N_VPWR_c_1827_n 0.00445602f $X=10.885 $Y=2.465 $X2=0
+ $Y2=0
cc_594 N_RESET_B_c_568_n N_VPWR_c_1813_n 0.00453497f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_595 N_RESET_B_c_571_n N_VPWR_c_1813_n 9.43083e-19 $X=7.685 $Y=2.23 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_574_n N_VPWR_c_1813_n 0.00896147f $X=10.885 $Y=2.465 $X2=0
+ $Y2=0
cc_597 N_RESET_B_M1016_g N_A_300_464#_c_1975_n 0.0119496f $X=3.655 $Y=0.615
+ $X2=0 $Y2=0
cc_598 N_RESET_B_c_568_n N_A_300_464#_c_1976_n 0.0195497f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_599 N_RESET_B_M1016_g N_A_300_464#_c_1976_n 0.0263571f $X=3.655 $Y=0.615
+ $X2=0 $Y2=0
cc_600 N_RESET_B_c_576_n N_A_300_464#_c_1976_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_601 N_RESET_B_c_582_n N_A_300_464#_c_1976_n 0.0228135f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_602 N_RESET_B_c_575_n N_A_300_464#_c_1984_n 0.0290302f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_603 N_RESET_B_c_576_n N_A_300_464#_c_1984_n 0.00388056f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_604 N_RESET_B_c_581_n N_A_300_464#_c_1984_n 0.00258186f $X=3.95 $Y=1.995
+ $X2=0 $Y2=0
cc_605 N_RESET_B_c_582_n N_A_300_464#_c_1984_n 0.00903824f $X=3.95 $Y=1.995
+ $X2=0 $Y2=0
cc_606 N_RESET_B_c_568_n N_A_300_464#_c_1985_n 0.0205728f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_607 N_RESET_B_c_576_n N_A_300_464#_c_1985_n 4.98701e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_RESET_B_c_582_n N_A_300_464#_c_1985_n 0.0168153f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_575_n N_A_300_464#_c_1978_n 0.00362547f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_610 N_RESET_B_c_575_n N_A_300_464#_c_1987_n 0.0179072f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_611 N_RESET_B_c_575_n N_A_300_464#_c_1988_n 0.0167929f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_612 N_RESET_B_c_575_n N_A_300_464#_c_1980_n 0.0094217f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_613 N_RESET_B_c_568_n N_A_300_464#_c_1991_n 0.00629514f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_614 N_RESET_B_M1016_g N_VGND_c_2148_n 0.0028678f $X=3.655 $Y=0.615 $X2=0
+ $Y2=0
cc_615 N_RESET_B_M1038_g N_VGND_c_2150_n 0.00390833f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_616 N_RESET_B_M1016_g N_VGND_c_2153_n 0.00478603f $X=3.655 $Y=0.615 $X2=0
+ $Y2=0
cc_617 N_RESET_B_c_561_n N_VGND_c_2158_n 0.0033127f $X=7.3 $Y=1.085 $X2=0 $Y2=0
cc_618 N_RESET_B_M1038_g N_VGND_c_2160_n 0.00460063f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_619 N_RESET_B_M1016_g N_VGND_c_2163_n 0.0044912f $X=3.655 $Y=0.615 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_561_n N_VGND_c_2163_n 0.00479212f $X=7.3 $Y=1.085 $X2=0 $Y2=0
cc_621 N_RESET_B_M1038_g N_VGND_c_2163_n 0.00906826f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_622 N_RESET_B_M1016_g N_noxref_24_c_2273_n 0.0129714f $X=3.655 $Y=0.615 $X2=0
+ $Y2=0
cc_623 N_CLK_M1008_g N_A_1034_368#_c_828_n 6.18148e-19 $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_624 N_CLK_c_772_n N_A_1034_368#_c_832_n 8.47673e-19 $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_625 N_CLK_c_772_n N_A_855_368#_c_1280_n 0.0485382f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_626 N_CLK_M1008_g N_A_855_368#_c_1280_n 0.0260223f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_627 N_CLK_c_785_n N_A_855_368#_c_1280_n 2.65039e-19 $X=4.475 $Y=1.425 $X2=0
+ $Y2=0
cc_628 N_CLK_M1008_g N_A_855_368#_c_1281_n 0.0220186f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_629 N_CLK_M1008_g N_A_855_368#_c_1292_n 8.21824e-19 $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_630 N_CLK_M1008_g N_A_855_368#_c_1336_n 0.0146908f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_631 N_CLK_c_785_n N_A_855_368#_c_1336_n 0.00556295f $X=4.475 $Y=1.425 $X2=0
+ $Y2=0
cc_632 N_CLK_c_774_n N_A_855_368#_c_1322_n 0.00395112f $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_633 N_CLK_c_785_n N_A_855_368#_c_1322_n 0.0139041f $X=4.475 $Y=1.425 $X2=0
+ $Y2=0
cc_634 N_CLK_c_772_n N_A_855_368#_c_1310_n 0.011706f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_635 N_CLK_c_785_n N_A_855_368#_c_1310_n 0.00277151f $X=4.475 $Y=1.425 $X2=0
+ $Y2=0
cc_636 N_CLK_M1008_g N_A_855_368#_c_1293_n 0.00330582f $X=4.665 $Y=0.74 $X2=0
+ $Y2=0
cc_637 N_CLK_c_785_n N_A_855_368#_c_1293_n 0.00311452f $X=4.475 $Y=1.425 $X2=0
+ $Y2=0
cc_638 N_CLK_c_775_n N_A_855_368#_c_1293_n 0.00246687f $X=4.195 $Y=1.385 $X2=0
+ $Y2=0
cc_639 N_CLK_c_772_n N_A_855_368#_c_1294_n 0.00439259f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_640 N_CLK_c_772_n N_A_855_368#_c_1312_n 0.00541631f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_641 N_CLK_c_774_n N_A_855_368#_c_1312_n 0.004824f $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_642 N_CLK_c_785_n N_A_855_368#_c_1312_n 0.0144756f $X=4.475 $Y=1.425 $X2=0
+ $Y2=0
cc_643 N_CLK_c_772_n N_A_855_368#_c_1295_n 0.00338092f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_644 N_CLK_c_785_n N_A_855_368#_c_1295_n 0.0249312f $X=4.475 $Y=1.425 $X2=0
+ $Y2=0
cc_645 N_CLK_c_772_n N_VPWR_c_1816_n 0.0172823f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_646 N_CLK_c_772_n N_VPWR_c_1823_n 0.00413917f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_647 N_CLK_c_772_n N_VPWR_c_1813_n 0.00403443f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_648 N_CLK_c_774_n N_A_300_464#_c_1976_n 3.52805e-19 $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_649 N_CLK_c_775_n N_A_300_464#_c_1976_n 0.0189245f $X=4.195 $Y=1.385 $X2=0
+ $Y2=0
cc_650 N_CLK_c_772_n N_A_300_464#_c_1984_n 0.0146064f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_651 N_CLK_c_772_n N_A_300_464#_c_1985_n 0.00160388f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_652 N_CLK_c_772_n N_A_300_464#_c_1991_n 0.0102085f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_653 N_CLK_M1008_g N_VGND_c_2148_n 0.00313842f $X=4.665 $Y=0.74 $X2=0 $Y2=0
cc_654 N_CLK_M1008_g N_VGND_c_2149_n 0.010966f $X=4.665 $Y=0.74 $X2=0 $Y2=0
cc_655 N_CLK_M1008_g N_VGND_c_2155_n 0.00383152f $X=4.665 $Y=0.74 $X2=0 $Y2=0
cc_656 N_CLK_M1008_g N_VGND_c_2163_n 0.00762539f $X=4.665 $Y=0.74 $X2=0 $Y2=0
cc_657 N_A_1034_368#_c_836_n N_A_1367_92#_M1033_d 0.00176461f $X=9.065 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_658 N_A_1034_368#_M1000_g N_A_1367_92#_M1027_g 0.0326305f $X=6.52 $Y=0.8
+ $X2=0 $Y2=0
cc_659 N_A_1034_368#_c_830_n N_A_1367_92#_M1027_g 0.00660604f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_660 N_A_1034_368#_c_834_n N_A_1367_92#_M1027_g 0.00274482f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_661 N_A_1034_368#_c_872_p N_A_1367_92#_M1027_g 0.0026982f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_662 N_A_1034_368#_c_824_n N_A_1367_92#_c_1039_n 0.0326305f $X=6.445 $Y=1.65
+ $X2=0 $Y2=0
cc_663 N_A_1034_368#_c_843_n N_A_1367_92#_c_1039_n 0.00102464f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_664 N_A_1034_368#_c_835_n N_A_1367_92#_c_1040_n 0.0520185f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_665 N_A_1034_368#_c_836_n N_A_1367_92#_c_1040_n 0.00353238f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_666 N_A_1034_368#_c_835_n N_A_1367_92#_c_1041_n 0.00761753f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_667 N_A_1034_368#_c_872_p N_A_1367_92#_c_1041_n 0.0103944f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_668 N_A_1034_368#_c_839_n N_A_1367_92#_c_1048_n 0.0139231f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_669 N_A_1034_368#_c_844_n N_A_1367_92#_c_1048_n 0.00323506f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_670 N_A_1034_368#_c_826_n N_A_1367_92#_c_1042_n 0.014712f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_671 N_A_1034_368#_c_827_n N_A_1367_92#_c_1042_n 0.00243289f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_672 N_A_1034_368#_c_836_n N_A_1367_92#_c_1042_n 0.0257761f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_673 N_A_1034_368#_c_838_n N_A_1367_92#_c_1042_n 0.0141828f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_674 N_A_1034_368#_c_841_n N_A_1367_92#_c_1042_n 5.79172e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_675 N_A_1034_368#_c_842_n N_A_1367_92#_c_1042_n 0.0131302f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_676 N_A_1034_368#_c_844_n N_A_1367_92#_c_1042_n 0.00313966f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_677 N_A_1034_368#_c_839_n N_A_1367_92#_c_1043_n 0.0197161f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_678 N_A_1034_368#_c_841_n N_A_1367_92#_c_1043_n 2.26254e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_679 N_A_1034_368#_c_842_n N_A_1367_92#_c_1043_n 0.0131446f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_680 N_A_1034_368#_c_844_n N_A_1367_92#_c_1043_n 0.00960948f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_681 N_A_1034_368#_c_826_n N_A_1233_118#_M1033_g 0.0286306f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_682 N_A_1034_368#_c_836_n N_A_1233_118#_M1033_g 0.0116373f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_683 N_A_1034_368#_c_827_n N_A_1233_118#_c_1147_n 0.0152066f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_684 N_A_1034_368#_c_839_n N_A_1233_118#_c_1147_n 4.45404e-19 $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_685 N_A_1034_368#_c_846_n N_A_1233_118#_c_1157_n 0.00187655f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_686 N_A_1034_368#_c_824_n N_A_1233_118#_c_1157_n 7.04121e-19 $X=6.445 $Y=1.65
+ $X2=0 $Y2=0
cc_687 N_A_1034_368#_M1000_g N_A_1233_118#_c_1148_n 0.0100665f $X=6.52 $Y=0.8
+ $X2=0 $Y2=0
cc_688 N_A_1034_368#_c_830_n N_A_1233_118#_c_1148_n 0.0118561f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_689 N_A_1034_368#_c_845_n N_A_1233_118#_c_1149_n 6.14864e-19 $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_690 N_A_1034_368#_c_846_n N_A_1233_118#_c_1149_n 3.40922e-19 $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_691 N_A_1034_368#_M1000_g N_A_1233_118#_c_1149_n 0.00685047f $X=6.52 $Y=0.8
+ $X2=0 $Y2=0
cc_692 N_A_1034_368#_c_824_n N_A_1233_118#_c_1154_n 4.6222e-19 $X=6.445 $Y=1.65
+ $X2=0 $Y2=0
cc_693 N_A_1034_368#_M1000_g N_A_1233_118#_c_1154_n 0.00668439f $X=6.52 $Y=0.8
+ $X2=0 $Y2=0
cc_694 N_A_1034_368#_c_830_n N_A_1233_118#_c_1154_n 0.0202257f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_695 N_A_1034_368#_c_872_p N_A_1233_118#_c_1154_n 0.00487041f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_696 N_A_1034_368#_c_829_n N_A_855_368#_c_1280_n 6.45062e-19 $X=5.535 $Y=1.545
+ $X2=0 $Y2=0
cc_697 N_A_1034_368#_c_832_n N_A_855_368#_c_1280_n 0.010981f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_698 N_A_1034_368#_c_840_n N_A_855_368#_c_1280_n 0.00906399f $X=5.385 $Y=1.13
+ $X2=0 $Y2=0
cc_699 N_A_1034_368#_c_828_n N_A_855_368#_c_1281_n 0.00742047f $X=5.315 $Y=0.515
+ $X2=0 $Y2=0
cc_700 N_A_1034_368#_c_829_n N_A_855_368#_c_1281_n 0.0010546f $X=5.535 $Y=1.545
+ $X2=0 $Y2=0
cc_701 N_A_1034_368#_c_831_n N_A_855_368#_c_1281_n 0.00466613f $X=5.62 $Y=0.34
+ $X2=0 $Y2=0
cc_702 N_A_1034_368#_c_840_n N_A_855_368#_c_1281_n 0.00334153f $X=5.385 $Y=1.13
+ $X2=0 $Y2=0
cc_703 N_A_1034_368#_c_829_n N_A_855_368#_c_1282_n 0.00667209f $X=5.535 $Y=1.545
+ $X2=0 $Y2=0
cc_704 N_A_1034_368#_c_832_n N_A_855_368#_c_1282_n 0.00218784f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_705 N_A_1034_368#_c_845_n N_A_855_368#_c_1283_n 0.0111395f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_706 N_A_1034_368#_c_846_n N_A_855_368#_c_1283_n 0.0129863f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_707 N_A_1034_368#_c_829_n N_A_855_368#_c_1283_n 0.00999835f $X=5.535 $Y=1.545
+ $X2=0 $Y2=0
cc_708 N_A_1034_368#_c_832_n N_A_855_368#_c_1283_n 0.0180665f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_709 N_A_1034_368#_c_833_n N_A_855_368#_c_1283_n 0.00967807f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_710 N_A_1034_368#_c_843_n N_A_855_368#_c_1283_n 0.0213708f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_711 N_A_1034_368#_c_833_n N_A_855_368#_c_1284_n 0.00459232f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_712 N_A_1034_368#_c_843_n N_A_855_368#_c_1284_n 0.0170495f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_713 N_A_1034_368#_c_846_n N_A_855_368#_c_1298_n 0.00899632f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_714 N_A_1034_368#_M1000_g N_A_855_368#_M1009_g 0.0222935f $X=6.52 $Y=0.8
+ $X2=0 $Y2=0
cc_715 N_A_1034_368#_c_828_n N_A_855_368#_M1009_g 0.00517237f $X=5.315 $Y=0.515
+ $X2=0 $Y2=0
cc_716 N_A_1034_368#_c_830_n N_A_855_368#_M1009_g 0.00680216f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_717 N_A_1034_368#_c_846_n N_A_855_368#_c_1300_n 0.00151278f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_718 N_A_1034_368#_c_846_n N_A_855_368#_c_1302_n 0.0132738f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_719 N_A_1034_368#_c_824_n N_A_855_368#_c_1302_n 9.41757e-19 $X=6.445 $Y=1.65
+ $X2=0 $Y2=0
cc_720 N_A_1034_368#_c_848_n N_A_855_368#_c_1304_n 0.00644632f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_721 N_A_1034_368#_c_848_n N_A_855_368#_M1004_g 0.0153501f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_722 N_A_1034_368#_c_839_n N_A_855_368#_M1004_g 0.00856179f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_723 N_A_1034_368#_c_848_n N_A_855_368#_c_1286_n 0.00418242f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_724 N_A_1034_368#_c_839_n N_A_855_368#_c_1286_n 0.0121351f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_725 N_A_1034_368#_c_852_n N_A_855_368#_c_1286_n 0.00479207f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_726 N_A_1034_368#_c_841_n N_A_855_368#_c_1287_n 0.019069f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_727 N_A_1034_368#_c_842_n N_A_855_368#_c_1287_n 0.00163879f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_728 N_A_1034_368#_c_844_n N_A_855_368#_c_1287_n 0.00141289f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_729 N_A_1034_368#_c_839_n N_A_855_368#_c_1288_n 0.00153175f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_730 N_A_1034_368#_c_836_n N_A_855_368#_M1007_g 0.00301232f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_731 N_A_1034_368#_c_838_n N_A_855_368#_M1007_g 0.00129859f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_732 N_A_1034_368#_c_841_n N_A_855_368#_M1007_g 0.00125371f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_733 N_A_1034_368#_c_829_n N_A_855_368#_c_1290_n 0.00513573f $X=5.535 $Y=1.545
+ $X2=0 $Y2=0
cc_734 N_A_1034_368#_c_841_n N_A_855_368#_c_1291_n 0.0194128f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_735 N_A_1034_368#_c_842_n N_A_855_368#_c_1291_n 3.65519e-19 $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_736 N_A_1034_368#_c_832_n N_A_855_368#_c_1310_n 0.00783925f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_737 N_A_1034_368#_c_829_n N_A_855_368#_c_1293_n 0.00543166f $X=5.535 $Y=1.545
+ $X2=0 $Y2=0
cc_738 N_A_1034_368#_c_840_n N_A_855_368#_c_1293_n 0.00229916f $X=5.385 $Y=1.13
+ $X2=0 $Y2=0
cc_739 N_A_1034_368#_c_832_n N_A_855_368#_c_1294_n 0.00785664f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_740 N_A_1034_368#_c_832_n N_A_855_368#_c_1312_n 0.00461694f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_741 N_A_1034_368#_c_829_n N_A_855_368#_c_1295_n 0.0187727f $X=5.535 $Y=1.545
+ $X2=0 $Y2=0
cc_742 N_A_1034_368#_c_832_n N_A_855_368#_c_1295_n 0.0158577f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_743 N_A_1034_368#_c_840_n N_A_855_368#_c_1295_n 0.0107724f $X=5.385 $Y=1.13
+ $X2=0 $Y2=0
cc_744 N_A_1034_368#_c_848_n N_A_1997_272#_c_1494_n 0.0218756f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_745 N_A_1034_368#_c_852_n N_A_1997_272#_c_1494_n 2.75032e-19 $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_746 N_A_1034_368#_c_848_n N_A_1997_272#_c_1495_n 0.0293409f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_747 N_A_1034_368#_c_836_n N_A_1745_74#_M1010_d 0.00630965f $X=9.065 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_748 N_A_1034_368#_c_838_n N_A_1745_74#_M1010_d 0.0113887f $X=9.15 $Y=0.94
+ $X2=-0.19 $Y2=-0.245
cc_749 N_A_1034_368#_c_839_n N_A_1745_74#_M1004_d 0.00749069f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_750 N_A_1034_368#_c_961_p N_A_1745_74#_M1004_d 0.0039098f $X=9.415 $Y=2.252
+ $X2=0 $Y2=0
cc_751 N_A_1034_368#_c_852_n N_A_1745_74#_M1004_d 0.00176657f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_752 N_A_1034_368#_c_848_n N_A_1745_74#_c_1616_n 0.0220662f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_753 N_A_1034_368#_c_961_p N_A_1745_74#_c_1616_n 0.0101735f $X=9.415 $Y=2.252
+ $X2=0 $Y2=0
cc_754 N_A_1034_368#_c_852_n N_A_1745_74#_c_1616_n 0.0386883f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_755 N_A_1034_368#_c_838_n N_A_1745_74#_c_1604_n 0.00768735f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_756 N_A_1034_368#_c_841_n N_A_1745_74#_c_1604_n 4.55554e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_757 N_A_1034_368#_c_842_n N_A_1745_74#_c_1604_n 0.0116456f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_758 N_A_1034_368#_c_839_n N_A_1745_74#_c_1605_n 0.0375442f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_759 N_A_1034_368#_c_848_n N_A_1745_74#_c_1618_n 0.00443076f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_760 N_A_1034_368#_c_852_n N_A_1745_74#_c_1618_n 0.0125258f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_761 N_A_1034_368#_c_848_n N_A_1745_74#_c_1619_n 9.16255e-19 $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_762 N_A_1034_368#_c_839_n N_A_1745_74#_c_1619_n 0.0141314f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_763 N_A_1034_368#_c_852_n N_A_1745_74#_c_1619_n 0.0111216f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_764 N_A_1034_368#_c_848_n N_A_1745_74#_c_1620_n 0.0062593f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_765 N_A_1034_368#_c_852_n N_A_1745_74#_c_1620_n 0.0202186f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_766 N_A_1034_368#_c_826_n N_A_1745_74#_c_1606_n 5.77109e-19 $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_767 N_A_1034_368#_c_836_n N_A_1745_74#_c_1606_n 0.00648023f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_768 N_A_1034_368#_c_838_n N_A_1745_74#_c_1606_n 0.0264512f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_769 N_A_1034_368#_c_841_n N_A_1745_74#_c_1606_n 2.06488e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_770 N_A_1034_368#_c_842_n N_A_1745_74#_c_1606_n 7.15367e-19 $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_771 N_A_1034_368#_c_841_n N_A_1745_74#_c_1607_n 6.39686e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_772 N_A_1034_368#_c_842_n N_A_1745_74#_c_1607_n 0.0144646f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_773 N_A_1034_368#_c_848_n N_VPWR_c_1825_n 0.00304676f $X=9.89 $Y=2.465 $X2=0
+ $Y2=0
cc_774 N_A_1034_368#_c_846_n N_VPWR_c_1813_n 9.49986e-19 $X=6.135 $Y=2.21 $X2=0
+ $Y2=0
cc_775 N_A_1034_368#_c_848_n N_VPWR_c_1813_n 0.00375875f $X=9.89 $Y=2.465 $X2=0
+ $Y2=0
cc_776 N_A_1034_368#_M1029_d N_A_300_464#_c_1984_n 0.00696197f $X=5.17 $Y=1.84
+ $X2=0 $Y2=0
cc_777 N_A_1034_368#_c_832_n N_A_300_464#_c_1984_n 0.0299967f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_778 N_A_1034_368#_c_833_n N_A_300_464#_c_1984_n 0.00299482f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_779 N_A_1034_368#_c_828_n N_A_300_464#_c_1977_n 0.0481284f $X=5.315 $Y=0.515
+ $X2=0 $Y2=0
cc_780 N_A_1034_368#_c_830_n N_A_300_464#_c_1977_n 0.012971f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_781 N_A_1034_368#_c_846_n N_A_300_464#_c_1986_n 0.00792141f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_782 N_A_1034_368#_c_832_n N_A_300_464#_c_1986_n 3.11389e-19 $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_783 N_A_1034_368#_c_824_n N_A_300_464#_c_1978_n 0.00319576f $X=6.445 $Y=1.65
+ $X2=0 $Y2=0
cc_784 N_A_1034_368#_M1000_g N_A_300_464#_c_1978_n 0.00628679f $X=6.52 $Y=0.8
+ $X2=0 $Y2=0
cc_785 N_A_1034_368#_c_833_n N_A_300_464#_c_1978_n 0.0171336f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_786 N_A_1034_368#_c_843_n N_A_300_464#_c_1978_n 0.00297767f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_787 N_A_1034_368#_c_829_n N_A_300_464#_c_1979_n 0.0130742f $X=5.535 $Y=1.545
+ $X2=0 $Y2=0
cc_788 N_A_1034_368#_c_833_n N_A_300_464#_c_1979_n 0.0140665f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_789 N_A_1034_368#_c_843_n N_A_300_464#_c_1979_n 3.69257e-19 $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_790 N_A_1034_368#_c_845_n N_A_300_464#_c_1987_n 0.00392277f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_791 N_A_1034_368#_c_846_n N_A_300_464#_c_1987_n 0.00875358f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_792 N_A_1034_368#_c_824_n N_A_300_464#_c_1987_n 0.00254238f $X=6.445 $Y=1.65
+ $X2=0 $Y2=0
cc_793 N_A_1034_368#_c_833_n N_A_300_464#_c_1987_n 0.00770757f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_794 N_A_1034_368#_c_845_n N_A_300_464#_c_1988_n 0.00121768f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_795 N_A_1034_368#_c_846_n N_A_300_464#_c_1988_n 0.00154832f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_796 N_A_1034_368#_c_832_n N_A_300_464#_c_1988_n 0.0117904f $X=5.62 $Y=1.71
+ $X2=0 $Y2=0
cc_797 N_A_1034_368#_c_833_n N_A_300_464#_c_1988_n 0.0168093f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_798 N_A_1034_368#_c_843_n N_A_300_464#_c_1988_n 0.00323248f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_799 N_A_1034_368#_c_845_n N_A_300_464#_c_1980_n 0.00549102f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_800 N_A_1034_368#_c_824_n N_A_300_464#_c_1980_n 0.0105431f $X=6.445 $Y=1.65
+ $X2=0 $Y2=0
cc_801 N_A_1034_368#_M1000_g N_A_300_464#_c_1980_n 0.00582859f $X=6.52 $Y=0.8
+ $X2=0 $Y2=0
cc_802 N_A_1034_368#_c_833_n N_A_300_464#_c_1980_n 0.0256508f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_803 N_A_1034_368#_c_843_n N_A_300_464#_c_1980_n 0.00265891f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_804 N_A_1034_368#_c_835_n N_VGND_M1019_d 0.0169732f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_805 N_A_1034_368#_c_862_n N_VGND_M1019_d 0.00350731f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_806 N_A_1034_368#_c_837_n N_VGND_M1019_d 0.00122695f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_807 N_A_1034_368#_c_828_n N_VGND_c_2149_n 0.0237343f $X=5.315 $Y=0.515 $X2=0
+ $Y2=0
cc_808 N_A_1034_368#_c_831_n N_VGND_c_2149_n 0.0130228f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_809 N_A_1034_368#_c_830_n N_VGND_c_2158_n 0.10396f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_810 N_A_1034_368#_c_831_n N_VGND_c_2158_n 0.0336049f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_811 N_A_1034_368#_c_835_n N_VGND_c_2158_n 0.00402072f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_812 N_A_1034_368#_c_826_n N_VGND_c_2159_n 0.00278271f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_813 N_A_1034_368#_c_835_n N_VGND_c_2159_n 0.00335833f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_814 N_A_1034_368#_c_836_n N_VGND_c_2159_n 0.0734255f $X=9.065 $Y=0.34 $X2=0
+ $Y2=0
cc_815 N_A_1034_368#_c_837_n N_VGND_c_2159_n 0.0118998f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_816 N_A_1034_368#_c_826_n N_VGND_c_2163_n 0.00358525f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_817 N_A_1034_368#_c_830_n N_VGND_c_2163_n 0.0603123f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_818 N_A_1034_368#_c_831_n N_VGND_c_2163_n 0.0181581f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_819 N_A_1034_368#_c_835_n N_VGND_c_2163_n 0.0128826f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_820 N_A_1034_368#_c_836_n N_VGND_c_2163_n 0.0415191f $X=9.065 $Y=0.34 $X2=0
+ $Y2=0
cc_821 N_A_1034_368#_c_837_n N_VGND_c_2163_n 0.00655543f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_822 N_A_1034_368#_c_830_n N_VGND_c_2165_n 0.0118145f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_823 N_A_1034_368#_c_835_n N_VGND_c_2165_n 0.0246013f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_824 N_A_1034_368#_c_837_n N_VGND_c_2165_n 0.0135793f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_825 N_A_1034_368#_c_872_p A_1397_118# 0.00355812f $X=7.22 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_826 N_A_1367_92#_c_1040_n N_A_1233_118#_M1033_g 0.0106637f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_827 N_A_1367_92#_c_1042_n N_A_1233_118#_M1033_g 0.0114957f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_828 N_A_1367_92#_c_1043_n N_A_1233_118#_M1033_g 9.26224e-19 $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_829 N_A_1367_92#_c_1042_n N_A_1233_118#_c_1147_n 0.00716915f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_830 N_A_1367_92#_c_1043_n N_A_1233_118#_c_1147_n 0.0102608f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_831 N_A_1367_92#_c_1048_n N_A_1233_118#_c_1156_n 0.00282141f $X=8.865
+ $Y=1.855 $X2=0 $Y2=0
cc_832 N_A_1367_92#_c_1049_n N_A_1233_118#_c_1156_n 0.0109404f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_833 N_A_1367_92#_c_1043_n N_A_1233_118#_c_1156_n 0.00260822f $X=8.865
+ $Y=1.715 $X2=0 $Y2=0
cc_834 N_A_1367_92#_M1027_g N_A_1233_118#_c_1148_n 0.00505673f $X=6.91 $Y=0.8
+ $X2=0 $Y2=0
cc_835 N_A_1367_92#_c_1041_n N_A_1233_118#_c_1148_n 0.00930726f $X=7.325
+ $Y=1.005 $X2=0 $Y2=0
cc_836 N_A_1367_92#_M1027_g N_A_1233_118#_c_1149_n 0.00779885f $X=6.91 $Y=0.8
+ $X2=0 $Y2=0
cc_837 N_A_1367_92#_c_1044_n N_A_1233_118#_c_1149_n 0.00991263f $X=7.06 $Y=2.14
+ $X2=0 $Y2=0
cc_838 N_A_1367_92#_c_1045_n N_A_1233_118#_c_1149_n 9.97148e-19 $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_839 N_A_1367_92#_c_1038_n N_A_1233_118#_c_1149_n 0.0517809f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_840 N_A_1367_92#_c_1039_n N_A_1233_118#_c_1149_n 0.00941718f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_841 N_A_1367_92#_c_1041_n N_A_1233_118#_c_1149_n 0.00480628f $X=7.325
+ $Y=1.005 $X2=0 $Y2=0
cc_842 N_A_1367_92#_c_1045_n N_A_1233_118#_c_1168_n 0.0116684f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_843 N_A_1367_92#_c_1038_n N_A_1233_118#_c_1168_n 0.0034045f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_844 N_A_1367_92#_c_1039_n N_A_1233_118#_c_1168_n 0.00356794f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_845 N_A_1367_92#_c_1044_n N_A_1233_118#_c_1150_n 0.00330246f $X=7.06 $Y=2.14
+ $X2=0 $Y2=0
cc_846 N_A_1367_92#_c_1045_n N_A_1233_118#_c_1150_n 0.00151519f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_847 N_A_1367_92#_c_1038_n N_A_1233_118#_c_1150_n 0.0170101f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_848 N_A_1367_92#_c_1039_n N_A_1233_118#_c_1150_n 0.00147646f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_849 N_A_1367_92#_c_1038_n N_A_1233_118#_c_1151_n 0.0271019f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_850 N_A_1367_92#_c_1039_n N_A_1233_118#_c_1151_n 7.33487e-19 $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_851 N_A_1367_92#_c_1040_n N_A_1233_118#_c_1151_n 0.0133652f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_852 N_A_1367_92#_c_1040_n N_A_1233_118#_c_1152_n 0.0454545f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_853 N_A_1367_92#_c_1042_n N_A_1233_118#_c_1152_n 0.00357705f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_854 N_A_1367_92#_c_1043_n N_A_1233_118#_c_1152_n 0.0123924f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_855 N_A_1367_92#_c_1040_n N_A_1233_118#_c_1153_n 0.00365093f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_856 N_A_1367_92#_c_1042_n N_A_1233_118#_c_1153_n 4.74815e-19 $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_857 N_A_1367_92#_c_1043_n N_A_1233_118#_c_1153_n 0.00153128f $X=8.865
+ $Y=1.715 $X2=0 $Y2=0
cc_858 N_A_1367_92#_M1027_g N_A_1233_118#_c_1154_n 0.00108182f $X=6.91 $Y=0.8
+ $X2=0 $Y2=0
cc_859 N_A_1367_92#_c_1045_n N_A_1233_118#_c_1161_n 0.00554019f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_860 N_A_1367_92#_c_1045_n N_A_855_368#_c_1300_n 0.00284772f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_861 N_A_1367_92#_c_1045_n N_A_855_368#_c_1302_n 0.0278287f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_862 N_A_1367_92#_c_1045_n N_A_855_368#_c_1303_n 0.0095327f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_863 N_A_1367_92#_c_1049_n N_A_855_368#_c_1303_n 0.00408637f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_864 N_A_1367_92#_c_1048_n N_A_855_368#_M1004_g 0.0075382f $X=8.865 $Y=1.855
+ $X2=0 $Y2=0
cc_865 N_A_1367_92#_c_1043_n N_A_855_368#_M1004_g 4.14175e-19 $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_866 N_A_1367_92#_c_1043_n N_A_855_368#_c_1287_n 0.00134852f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_867 N_A_1367_92#_c_1042_n N_A_1745_74#_M1010_d 0.00295216f $X=8.435 $Y=0.81
+ $X2=-0.19 $Y2=-0.245
cc_868 N_A_1367_92#_c_1049_n N_A_1745_74#_c_1616_n 0.0117842f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_869 N_A_1367_92#_c_1045_n N_VPWR_c_1817_n 0.00454716f $X=7.06 $Y=2.23 $X2=0
+ $Y2=0
cc_870 N_A_1367_92#_c_1048_n N_VPWR_c_1819_n 0.0728f $X=8.865 $Y=1.855 $X2=0
+ $Y2=0
cc_871 N_A_1367_92#_c_1042_n N_VPWR_c_1819_n 0.00559467f $X=8.435 $Y=0.81 $X2=0
+ $Y2=0
cc_872 N_A_1367_92#_c_1049_n N_VPWR_c_1825_n 0.00629779f $X=8.92 $Y=1.88 $X2=0
+ $Y2=0
cc_873 N_A_1367_92#_c_1045_n N_VPWR_c_1813_n 9.43083e-19 $X=7.06 $Y=2.23 $X2=0
+ $Y2=0
cc_874 N_A_1367_92#_c_1049_n N_VPWR_c_1813_n 0.00766223f $X=8.92 $Y=1.88 $X2=0
+ $Y2=0
cc_875 N_A_1367_92#_M1027_g N_A_300_464#_c_1980_n 3.2774e-19 $X=6.91 $Y=0.8
+ $X2=0 $Y2=0
cc_876 N_A_1367_92#_c_1039_n N_A_300_464#_c_1980_n 2.3169e-19 $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_877 N_A_1367_92#_c_1040_n N_VGND_M1019_d 0.00718336f $X=8.27 $Y=1.005 $X2=0
+ $Y2=0
cc_878 N_A_1367_92#_c_1041_n A_1397_118# 0.00206764f $X=7.325 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_879 N_A_1233_118#_c_1157_n N_A_855_368#_c_1298_n 0.00396944f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_880 N_A_1233_118#_c_1154_n N_A_855_368#_M1009_g 0.00579532f $X=6.305 $Y=0.81
+ $X2=0 $Y2=0
cc_881 N_A_1233_118#_c_1157_n N_A_855_368#_c_1302_n 0.00984149f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_882 N_A_1233_118#_c_1149_n N_A_855_368#_c_1302_n 0.00327177f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_883 N_A_1233_118#_c_1161_n N_A_855_368#_c_1302_n 0.00504398f $X=6.795
+ $Y=2.522 $X2=0 $Y2=0
cc_884 N_A_1233_118#_c_1156_n N_A_855_368#_c_1303_n 0.0102036f $X=8.695 $Y=1.66
+ $X2=0 $Y2=0
cc_885 N_A_1233_118#_c_1168_n N_A_855_368#_c_1303_n 0.003989f $X=7.495 $Y=2.405
+ $X2=0 $Y2=0
cc_886 N_A_1233_118#_c_1150_n N_A_855_368#_c_1303_n 0.00777265f $X=7.58 $Y=2.32
+ $X2=0 $Y2=0
cc_887 N_A_1233_118#_c_1161_n N_A_855_368#_c_1303_n 0.00119096f $X=6.795
+ $Y=2.522 $X2=0 $Y2=0
cc_888 N_A_1233_118#_c_1156_n N_A_855_368#_c_1304_n 0.00230914f $X=8.695 $Y=1.66
+ $X2=0 $Y2=0
cc_889 N_A_1233_118#_c_1156_n N_A_855_368#_M1004_g 0.00557664f $X=8.695 $Y=1.66
+ $X2=0 $Y2=0
cc_890 N_A_1233_118#_c_1147_n N_A_855_368#_c_1287_n 0.00717177f $X=8.605 $Y=1.52
+ $X2=0 $Y2=0
cc_891 N_A_1233_118#_c_1168_n N_VPWR_M1002_d 0.00772988f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_892 N_A_1233_118#_c_1150_n N_VPWR_M1002_d 7.78169e-19 $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_893 N_A_1233_118#_c_1168_n N_VPWR_c_1817_n 0.0222224f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_894 N_A_1233_118#_c_1150_n N_VPWR_c_1817_n 0.00949227f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_895 N_A_1233_118#_c_1161_n N_VPWR_c_1817_n 0.00341149f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_896 N_A_1233_118#_c_1150_n N_VPWR_c_1818_n 0.00714098f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_897 N_A_1233_118#_c_1147_n N_VPWR_c_1819_n 0.00460268f $X=8.605 $Y=1.52 $X2=0
+ $Y2=0
cc_898 N_A_1233_118#_c_1156_n N_VPWR_c_1819_n 0.00728995f $X=8.695 $Y=1.66 $X2=0
+ $Y2=0
cc_899 N_A_1233_118#_c_1150_n N_VPWR_c_1819_n 0.0222061f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_900 N_A_1233_118#_c_1157_n N_VPWR_c_1831_n 0.00833207f $X=6.71 $Y=2.555 $X2=0
+ $Y2=0
cc_901 N_A_1233_118#_c_1161_n N_VPWR_c_1831_n 0.00291643f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_902 N_A_1233_118#_c_1156_n N_VPWR_c_1813_n 9.39239e-19 $X=8.695 $Y=1.66 $X2=0
+ $Y2=0
cc_903 N_A_1233_118#_c_1157_n N_VPWR_c_1813_n 0.0118132f $X=6.71 $Y=2.555 $X2=0
+ $Y2=0
cc_904 N_A_1233_118#_c_1168_n N_VPWR_c_1813_n 0.0104334f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_905 N_A_1233_118#_c_1150_n N_VPWR_c_1813_n 0.0154819f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_906 N_A_1233_118#_c_1161_n N_VPWR_c_1813_n 0.00457064f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_907 N_A_1233_118#_c_1154_n N_A_300_464#_c_1977_n 0.0162775f $X=6.305 $Y=0.81
+ $X2=0 $Y2=0
cc_908 N_A_1233_118#_c_1157_n N_A_300_464#_c_1986_n 0.0136661f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_909 N_A_1233_118#_c_1149_n N_A_300_464#_c_1986_n 0.00242728f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_910 N_A_1233_118#_c_1161_n N_A_300_464#_c_1986_n 0.00169407f $X=6.795
+ $Y=2.522 $X2=0 $Y2=0
cc_911 N_A_1233_118#_c_1148_n N_A_300_464#_c_1978_n 0.00533227f $X=6.71 $Y=0.945
+ $X2=0 $Y2=0
cc_912 N_A_1233_118#_c_1149_n N_A_300_464#_c_1978_n 0.0135848f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_913 N_A_1233_118#_c_1154_n N_A_300_464#_c_1978_n 0.0271808f $X=6.305 $Y=0.81
+ $X2=0 $Y2=0
cc_914 N_A_1233_118#_c_1157_n N_A_300_464#_c_1987_n 0.0207396f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_915 N_A_1233_118#_c_1149_n N_A_300_464#_c_1987_n 0.0135339f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_916 N_A_1233_118#_c_1149_n N_A_300_464#_c_1980_n 0.049001f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_917 N_A_1233_118#_c_1168_n A_1343_461# 6.70978e-19 $X=7.495 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_918 N_A_1233_118#_c_1161_n A_1343_461# 0.00461414f $X=6.795 $Y=2.522
+ $X2=-0.19 $Y2=-0.245
cc_919 N_A_1233_118#_M1033_g N_VGND_c_2159_n 0.00278271f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_920 N_A_1233_118#_M1033_g N_VGND_c_2163_n 0.00358525f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_921 N_A_1233_118#_M1033_g N_VGND_c_2165_n 0.00111149f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_922 N_A_1233_118#_c_1148_n A_1319_118# 0.00209187f $X=6.71 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_923 N_A_855_368#_c_1288_n N_A_1997_272#_M1005_g 0.0100846f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_924 N_A_855_368#_M1007_g N_A_1997_272#_M1005_g 0.0520068f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_925 N_A_855_368#_c_1288_n N_A_1997_272#_c_1483_n 0.019486f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_926 N_A_855_368#_c_1288_n N_A_1997_272#_c_1490_n 6.49074e-19 $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_927 N_A_855_368#_c_1304_n N_A_1745_74#_c_1616_n 0.00244716f $X=9.145 $Y=2.9
+ $X2=0 $Y2=0
cc_928 N_A_855_368#_M1004_g N_A_1745_74#_c_1616_n 0.00467021f $X=9.145 $Y=2.235
+ $X2=0 $Y2=0
cc_929 N_A_855_368#_M1007_g N_A_1745_74#_c_1604_n 0.00653104f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_930 N_A_855_368#_c_1291_n N_A_1745_74#_c_1604_n 0.00549286f $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_931 N_A_855_368#_c_1286_n N_A_1745_74#_c_1605_n 0.0090777f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_932 N_A_855_368#_c_1288_n N_A_1745_74#_c_1605_n 0.00911046f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_933 N_A_855_368#_c_1286_n N_A_1745_74#_c_1618_n 2.60059e-19 $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_934 N_A_855_368#_c_1291_n N_A_1745_74#_c_1618_n 3.58986e-19 $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_935 N_A_855_368#_M1007_g N_A_1745_74#_c_1606_n 0.00822927f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_936 N_A_855_368#_c_1288_n N_A_1745_74#_c_1607_n 0.00212136f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_937 N_A_855_368#_c_1291_n N_A_1745_74#_c_1607_n 3.68292e-19 $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_938 N_A_855_368#_c_1288_n N_A_1745_74#_c_1609_n 0.00241471f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_939 N_A_855_368#_c_1291_n N_A_1745_74#_c_1609_n 0.00651625f $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_940 N_A_855_368#_c_1310_n N_VPWR_M1022_d 0.0023266f $X=4.81 $Y=1.905 $X2=0
+ $Y2=0
cc_941 N_A_855_368#_c_1280_n N_VPWR_c_1816_n 0.00888208f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_942 N_A_855_368#_c_1283_n N_VPWR_c_1816_n 0.0017658f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_943 N_A_855_368#_c_1299_n N_VPWR_c_1816_n 0.00232909f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_944 N_A_855_368#_c_1300_n N_VPWR_c_1817_n 0.00612345f $X=6.64 $Y=2.89 $X2=0
+ $Y2=0
cc_945 N_A_855_368#_c_1303_n N_VPWR_c_1817_n 0.025635f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_946 N_A_855_368#_c_1303_n N_VPWR_c_1818_n 0.0260958f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_947 N_A_855_368#_c_1303_n N_VPWR_c_1819_n 0.0170937f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_948 N_A_855_368#_c_1304_n N_VPWR_c_1819_n 0.00527525f $X=9.145 $Y=2.9 $X2=0
+ $Y2=0
cc_949 N_A_855_368#_c_1303_n N_VPWR_c_1825_n 0.0217861f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_950 N_A_855_368#_c_1280_n N_VPWR_c_1831_n 0.00413917f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_951 N_A_855_368#_c_1299_n N_VPWR_c_1831_n 0.0512154f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_952 N_A_855_368#_c_1280_n N_VPWR_c_1813_n 0.00399275f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_953 N_A_855_368#_c_1298_n N_VPWR_c_1813_n 0.0252643f $X=6.55 $Y=3.15 $X2=0
+ $Y2=0
cc_954 N_A_855_368#_c_1299_n N_VPWR_c_1813_n 0.00693725f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_955 N_A_855_368#_c_1303_n N_VPWR_c_1813_n 0.0749028f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_956 N_A_855_368#_c_1309_n N_VPWR_c_1813_n 0.00503906f $X=6.64 $Y=3.15 $X2=0
+ $Y2=0
cc_957 N_A_855_368#_M1022_s N_A_300_464#_c_1984_n 0.0082239f $X=4.275 $Y=1.84
+ $X2=0 $Y2=0
cc_958 N_A_855_368#_c_1280_n N_A_300_464#_c_1984_n 0.0126398f $X=5.095 $Y=1.765
+ $X2=0 $Y2=0
cc_959 N_A_855_368#_c_1283_n N_A_300_464#_c_1984_n 0.0133f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_960 N_A_855_368#_c_1298_n N_A_300_464#_c_1984_n 0.00106149f $X=6.55 $Y=3.15
+ $X2=0 $Y2=0
cc_961 N_A_855_368#_c_1310_n N_A_300_464#_c_1984_n 0.00793285f $X=4.81 $Y=1.905
+ $X2=0 $Y2=0
cc_962 N_A_855_368#_c_1312_n N_A_300_464#_c_1984_n 0.013838f $X=4.46 $Y=1.905
+ $X2=0 $Y2=0
cc_963 N_A_855_368#_c_1281_n N_A_300_464#_c_1977_n 6.79826e-19 $X=5.1 $Y=1.185
+ $X2=0 $Y2=0
cc_964 N_A_855_368#_c_1284_n N_A_300_464#_c_1977_n 0.00375217f $X=6.015 $Y=1.26
+ $X2=0 $Y2=0
cc_965 N_A_855_368#_M1009_g N_A_300_464#_c_1977_n 0.00691426f $X=6.09 $Y=0.8
+ $X2=0 $Y2=0
cc_966 N_A_855_368#_c_1283_n N_A_300_464#_c_1986_n 0.00814963f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_967 N_A_855_368#_c_1298_n N_A_300_464#_c_1986_n 0.00469098f $X=6.55 $Y=3.15
+ $X2=0 $Y2=0
cc_968 N_A_855_368#_c_1302_n N_A_300_464#_c_1986_n 4.63022e-19 $X=6.64 $Y=2.8
+ $X2=0 $Y2=0
cc_969 N_A_855_368#_c_1284_n N_A_300_464#_c_1978_n 0.0128725f $X=6.015 $Y=1.26
+ $X2=0 $Y2=0
cc_970 N_A_855_368#_c_1284_n N_A_300_464#_c_1979_n 0.00586816f $X=6.015 $Y=1.26
+ $X2=0 $Y2=0
cc_971 N_A_855_368#_c_1302_n N_A_300_464#_c_1987_n 3.77807e-19 $X=6.64 $Y=2.8
+ $X2=0 $Y2=0
cc_972 N_A_855_368#_c_1283_n N_A_300_464#_c_1988_n 0.00128765f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_973 N_A_855_368#_c_1283_n N_A_300_464#_c_1980_n 0.00248092f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_974 N_A_855_368#_c_1336_n N_VGND_M1008_d 0.00247461f $X=4.81 $Y=1.005 $X2=0
+ $Y2=0
cc_975 N_A_855_368#_c_1293_n N_VGND_M1008_d 2.0961e-19 $X=4.895 $Y=1.3 $X2=0
+ $Y2=0
cc_976 N_A_855_368#_c_1292_n N_VGND_c_2148_n 0.0153062f $X=4.45 $Y=0.515 $X2=0
+ $Y2=0
cc_977 N_A_855_368#_c_1281_n N_VGND_c_2149_n 0.00247266f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_978 N_A_855_368#_c_1292_n N_VGND_c_2149_n 0.0144259f $X=4.45 $Y=0.515 $X2=0
+ $Y2=0
cc_979 N_A_855_368#_c_1336_n N_VGND_c_2149_n 0.016164f $X=4.81 $Y=1.005 $X2=0
+ $Y2=0
cc_980 N_A_855_368#_M1007_g N_VGND_c_2150_n 0.0018065f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_981 N_A_855_368#_c_1292_n N_VGND_c_2155_n 0.00749631f $X=4.45 $Y=0.515 $X2=0
+ $Y2=0
cc_982 N_A_855_368#_c_1281_n N_VGND_c_2158_n 0.00430908f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_983 N_A_855_368#_M1007_g N_VGND_c_2159_n 0.00411612f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_984 N_A_855_368#_c_1281_n N_VGND_c_2163_n 0.00820937f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_985 N_A_855_368#_M1007_g N_VGND_c_2163_n 0.00752295f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_986 N_A_855_368#_c_1292_n N_VGND_c_2163_n 0.0062048f $X=4.45 $Y=0.515 $X2=0
+ $Y2=0
cc_987 N_A_1997_272#_c_1485_n N_A_1745_74#_M1028_g 0.00755075f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_988 N_A_1997_272#_c_1488_n N_A_1745_74#_M1028_g 0.00686241f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_989 N_A_1997_272#_c_1489_n N_A_1745_74#_M1028_g 3.28981e-19 $X=11.65 $Y=1.445
+ $X2=0 $Y2=0
cc_990 N_A_1997_272#_c_1486_n N_A_1745_74#_c_1600_n 0.0096742f $X=11.565 $Y=1.53
+ $X2=0 $Y2=0
cc_991 N_A_1997_272#_c_1491_n N_A_1745_74#_c_1600_n 0.012401f $X=11.127 $Y=2.52
+ $X2=0 $Y2=0
cc_992 N_A_1997_272#_c_1492_n N_A_1745_74#_c_1600_n 0.00480843f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_993 N_A_1997_272#_c_1491_n N_A_1745_74#_c_1611_n 0.00856137f $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_994 N_A_1997_272#_c_1496_n N_A_1745_74#_c_1612_n 0.00688539f $X=11.11 $Y=2.75
+ $X2=0 $Y2=0
cc_995 N_A_1997_272#_c_1491_n N_A_1745_74#_c_1612_n 0.00314773f $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_996 N_A_1997_272#_c_1486_n N_A_1745_74#_c_1601_n 0.00243079f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_997 N_A_1997_272#_c_1487_n N_A_1745_74#_c_1601_n 0.00158858f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_998 N_A_1997_272#_c_1489_n N_A_1745_74#_c_1601_n 0.0150077f $X=11.65 $Y=1.445
+ $X2=0 $Y2=0
cc_999 N_A_1997_272#_c_1484_n N_A_1745_74#_c_1602_n 0.00191851f $X=11.14 $Y=1.53
+ $X2=0 $Y2=0
cc_1000 N_A_1997_272#_c_1487_n N_A_1745_74#_c_1602_n 0.00173828f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1001 N_A_1997_272#_c_1488_n N_A_1745_74#_c_1602_n 0.00908089f $X=11.34
+ $Y=0.84 $X2=0 $Y2=0
cc_1002 N_A_1997_272#_c_1489_n N_A_1745_74#_c_1602_n 0.00419353f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1003 N_A_1997_272#_c_1492_n N_A_1745_74#_c_1602_n 0.00279652f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_1004 N_A_1997_272#_c_1486_n N_A_1745_74#_c_1613_n 0.00200907f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1005 N_A_1997_272#_c_1491_n N_A_1745_74#_c_1613_n 2.62811e-19 $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1006 N_A_1997_272#_c_1491_n N_A_1745_74#_c_1614_n 4.34489e-19 $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1007 N_A_1997_272#_c_1485_n N_A_1745_74#_M1031_g 0.00345625f $X=11.175
+ $Y=0.58 $X2=0 $Y2=0
cc_1008 N_A_1997_272#_c_1487_n N_A_1745_74#_M1031_g 0.00399686f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1009 N_A_1997_272#_c_1489_n N_A_1745_74#_M1031_g 0.00292154f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1010 N_A_1997_272#_c_1486_n N_A_1745_74#_c_1615_n 0.00270233f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1011 N_A_1997_272#_c_1491_n N_A_1745_74#_c_1615_n 0.00843513f $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1012 N_A_1997_272#_c_1495_n N_A_1745_74#_c_1616_n 0.00953641f $X=10.31
+ $Y=2.465 $X2=0 $Y2=0
cc_1013 N_A_1997_272#_M1005_g N_A_1745_74#_c_1605_n 5.63627e-19 $X=10.145
+ $Y=0.58 $X2=0 $Y2=0
cc_1014 N_A_1997_272#_c_1483_n N_A_1745_74#_c_1605_n 0.00475655f $X=10.31
+ $Y=1.84 $X2=0 $Y2=0
cc_1015 N_A_1997_272#_c_1490_n N_A_1745_74#_c_1605_n 0.0105779f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1016 N_A_1997_272#_c_1483_n N_A_1745_74#_c_1618_n 0.0112071f $X=10.31 $Y=1.84
+ $X2=0 $Y2=0
cc_1017 N_A_1997_272#_c_1494_n N_A_1745_74#_c_1618_n 0.00484392f $X=10.31
+ $Y=2.375 $X2=0 $Y2=0
cc_1018 N_A_1997_272#_c_1490_n N_A_1745_74#_c_1618_n 0.0232183f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1019 N_A_1997_272#_c_1494_n N_A_1745_74#_c_1620_n 0.011498f $X=10.31 $Y=2.375
+ $X2=0 $Y2=0
cc_1020 N_A_1997_272#_c_1495_n N_A_1745_74#_c_1620_n 0.00503711f $X=10.31
+ $Y=2.465 $X2=0 $Y2=0
cc_1021 N_A_1997_272#_M1005_g N_A_1745_74#_c_1606_n 0.00279105f $X=10.145
+ $Y=0.58 $X2=0 $Y2=0
cc_1022 N_A_1997_272#_c_1484_n N_A_1745_74#_c_1608_n 0.00534862f $X=11.14
+ $Y=1.53 $X2=0 $Y2=0
cc_1023 N_A_1997_272#_c_1486_n N_A_1745_74#_c_1608_n 0.0057529f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1024 N_A_1997_272#_c_1487_n N_A_1745_74#_c_1608_n 0.00391205f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1025 N_A_1997_272#_c_1489_n N_A_1745_74#_c_1608_n 0.0139087f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1026 N_A_1997_272#_c_1492_n N_A_1745_74#_c_1608_n 0.0134734f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_1027 N_A_1997_272#_M1005_g N_A_1745_74#_c_1609_n 0.0145056f $X=10.145 $Y=0.58
+ $X2=0 $Y2=0
cc_1028 N_A_1997_272#_c_1483_n N_A_1745_74#_c_1609_n 0.00481612f $X=10.31
+ $Y=1.84 $X2=0 $Y2=0
cc_1029 N_A_1997_272#_c_1484_n N_A_1745_74#_c_1609_n 0.0525955f $X=11.14 $Y=1.53
+ $X2=0 $Y2=0
cc_1030 N_A_1997_272#_c_1488_n N_A_1745_74#_c_1609_n 0.0263803f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_1031 N_A_1997_272#_c_1490_n N_A_1745_74#_c_1609_n 0.023139f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1032 N_A_1997_272#_c_1486_n N_A_2399_424#_c_1767_n 9.19806e-19 $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1033 N_A_1997_272#_c_1489_n N_A_2399_424#_c_1767_n 4.60428e-19 $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1034 N_A_1997_272#_c_1487_n N_A_2399_424#_c_1768_n 0.00457908f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1035 N_A_1997_272#_c_1489_n N_A_2399_424#_c_1768_n 0.0171651f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1036 N_A_1997_272#_c_1486_n N_A_2399_424#_c_1770_n 0.00962353f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1037 N_A_1997_272#_c_1489_n N_A_2399_424#_c_1770_n 0.00719431f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1038 N_A_1997_272#_c_1495_n N_VPWR_c_1820_n 0.00624782f $X=10.31 $Y=2.465
+ $X2=0 $Y2=0
cc_1039 N_A_1997_272#_c_1496_n N_VPWR_c_1820_n 0.0299967f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1040 N_A_1997_272#_c_1486_n N_VPWR_c_1821_n 0.0110039f $X=11.565 $Y=1.53
+ $X2=0 $Y2=0
cc_1041 N_A_1997_272#_c_1491_n N_VPWR_c_1821_n 0.067513f $X=11.127 $Y=2.52 $X2=0
+ $Y2=0
cc_1042 N_A_1997_272#_c_1495_n N_VPWR_c_1825_n 0.00377777f $X=10.31 $Y=2.465
+ $X2=0 $Y2=0
cc_1043 N_A_1997_272#_c_1496_n N_VPWR_c_1827_n 0.015771f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1044 N_A_1997_272#_c_1495_n N_VPWR_c_1813_n 0.00662633f $X=10.31 $Y=2.465
+ $X2=0 $Y2=0
cc_1045 N_A_1997_272#_c_1496_n N_VPWR_c_1813_n 0.0130108f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1046 N_A_1997_272#_c_1487_n N_VGND_M1031_s 0.00480139f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1047 N_A_1997_272#_M1005_g N_VGND_c_2150_n 0.01204f $X=10.145 $Y=0.58 $X2=0
+ $Y2=0
cc_1048 N_A_1997_272#_c_1485_n N_VGND_c_2150_n 0.0142227f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1049 N_A_1997_272#_c_1488_n N_VGND_c_2150_n 0.00176365f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_1050 N_A_1997_272#_c_1485_n N_VGND_c_2151_n 0.0158614f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1051 N_A_1997_272#_c_1487_n N_VGND_c_2151_n 0.0143444f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1052 N_A_1997_272#_M1005_g N_VGND_c_2159_n 0.00383152f $X=10.145 $Y=0.58
+ $X2=0 $Y2=0
cc_1053 N_A_1997_272#_c_1485_n N_VGND_c_2160_n 0.0143883f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1054 N_A_1997_272#_c_1487_n N_VGND_c_2160_n 0.00329108f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1055 N_A_1997_272#_M1005_g N_VGND_c_2163_n 0.0075694f $X=10.145 $Y=0.58 $X2=0
+ $Y2=0
cc_1056 N_A_1997_272#_c_1485_n N_VGND_c_2163_n 0.0119301f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1057 N_A_1997_272#_c_1487_n N_VGND_c_2163_n 0.00670825f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1058 N_A_1745_74#_c_1601_n N_A_2399_424#_c_1767_n 0.00328297f $X=11.88
+ $Y=1.275 $X2=0 $Y2=0
cc_1059 N_A_1745_74#_c_1613_n N_A_2399_424#_c_1773_n 7.20279e-19 $X=11.83
+ $Y=1.915 $X2=0 $Y2=0
cc_1060 N_A_1745_74#_c_1614_n N_A_2399_424#_c_1773_n 0.0133065f $X=11.92
+ $Y=2.045 $X2=0 $Y2=0
cc_1061 N_A_1745_74#_M1031_g N_A_2399_424#_c_1768_n 0.0137683f $X=11.955
+ $Y=0.645 $X2=0 $Y2=0
cc_1062 N_A_1745_74#_c_1600_n N_A_2399_424#_c_1769_n 0.00247742f $X=11.32
+ $Y=1.84 $X2=0 $Y2=0
cc_1063 N_A_1745_74#_c_1613_n N_A_2399_424#_c_1769_n 0.00929958f $X=11.83
+ $Y=1.915 $X2=0 $Y2=0
cc_1064 N_A_1745_74#_c_1614_n N_A_2399_424#_c_1769_n 0.00208502f $X=11.92
+ $Y=2.045 $X2=0 $Y2=0
cc_1065 N_A_1745_74#_c_1600_n N_A_2399_424#_c_1770_n 0.00108268f $X=11.32
+ $Y=1.84 $X2=0 $Y2=0
cc_1066 N_A_1745_74#_c_1601_n N_A_2399_424#_c_1770_n 5.99943e-19 $X=11.88
+ $Y=1.275 $X2=0 $Y2=0
cc_1067 N_A_1745_74#_c_1616_n N_VPWR_c_1820_n 0.0266532f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1068 N_A_1745_74#_c_1620_n N_VPWR_c_1820_n 0.00216548f $X=10.23 $Y=2.55 $X2=0
+ $Y2=0
cc_1069 N_A_1745_74#_c_1611_n N_VPWR_c_1821_n 0.00344007f $X=11.335 $Y=2.375
+ $X2=0 $Y2=0
cc_1070 N_A_1745_74#_c_1612_n N_VPWR_c_1821_n 0.00777412f $X=11.335 $Y=2.465
+ $X2=0 $Y2=0
cc_1071 N_A_1745_74#_c_1613_n N_VPWR_c_1821_n 0.0100207f $X=11.83 $Y=1.915 $X2=0
+ $Y2=0
cc_1072 N_A_1745_74#_c_1614_n N_VPWR_c_1821_n 0.00892462f $X=11.92 $Y=2.045
+ $X2=0 $Y2=0
cc_1073 N_A_1745_74#_c_1614_n N_VPWR_c_1822_n 0.00463887f $X=11.92 $Y=2.045
+ $X2=0 $Y2=0
cc_1074 N_A_1745_74#_c_1616_n N_VPWR_c_1825_n 0.0274952f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1075 N_A_1745_74#_c_1612_n N_VPWR_c_1827_n 0.00405947f $X=11.335 $Y=2.465
+ $X2=0 $Y2=0
cc_1076 N_A_1745_74#_c_1614_n N_VPWR_c_1832_n 0.00445602f $X=11.92 $Y=2.045
+ $X2=0 $Y2=0
cc_1077 N_A_1745_74#_c_1612_n N_VPWR_c_1813_n 0.00767502f $X=11.335 $Y=2.465
+ $X2=0 $Y2=0
cc_1078 N_A_1745_74#_c_1614_n N_VPWR_c_1813_n 0.00862869f $X=11.92 $Y=2.045
+ $X2=0 $Y2=0
cc_1079 N_A_1745_74#_c_1616_n N_VPWR_c_1813_n 0.0335089f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1080 N_A_1745_74#_c_1616_n A_1993_508# 0.00423971f $X=10.145 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1081 N_A_1745_74#_c_1606_n N_VGND_c_2150_n 0.0159689f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1082 N_A_1745_74#_c_1609_n N_VGND_c_2150_n 0.0191133f $X=11.065 $Y=1.185
+ $X2=0 $Y2=0
cc_1083 N_A_1745_74#_M1028_g N_VGND_c_2151_n 0.00322527f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1084 N_A_1745_74#_c_1601_n N_VGND_c_2151_n 0.00195495f $X=11.88 $Y=1.275
+ $X2=0 $Y2=0
cc_1085 N_A_1745_74#_M1031_g N_VGND_c_2151_n 0.00927494f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1086 N_A_1745_74#_M1031_g N_VGND_c_2152_n 0.00296233f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1087 N_A_1745_74#_c_1606_n N_VGND_c_2159_n 0.0151251f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1088 N_A_1745_74#_M1028_g N_VGND_c_2160_n 0.00434272f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1089 N_A_1745_74#_M1031_g N_VGND_c_2161_n 0.00383152f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1090 N_A_1745_74#_M1028_g N_VGND_c_2163_n 0.00825669f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1091 N_A_1745_74#_M1031_g N_VGND_c_2163_n 0.00762539f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1092 N_A_1745_74#_c_1606_n N_VGND_c_2163_n 0.0125365f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1093 N_A_2399_424#_c_1773_n N_VPWR_c_1821_n 0.0345631f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1094 N_A_2399_424#_c_1771_n N_VPWR_c_1822_n 0.0215785f $X=12.93 $Y=1.765
+ $X2=0 $Y2=0
cc_1095 N_A_2399_424#_c_1767_n N_VPWR_c_1822_n 0.00731242f $X=12.84 $Y=1.465
+ $X2=0 $Y2=0
cc_1096 N_A_2399_424#_c_1793_p N_VPWR_c_1822_n 0.0253438f $X=12.745 $Y=1.465
+ $X2=0 $Y2=0
cc_1097 N_A_2399_424#_c_1769_n N_VPWR_c_1822_n 0.0776081f $X=12.145 $Y=2.1 $X2=0
+ $Y2=0
cc_1098 N_A_2399_424#_c_1773_n N_VPWR_c_1832_n 0.0145938f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1099 N_A_2399_424#_c_1771_n N_VPWR_c_1833_n 0.00413917f $X=12.93 $Y=1.765
+ $X2=0 $Y2=0
cc_1100 N_A_2399_424#_c_1771_n N_VPWR_c_1813_n 0.00821237f $X=12.93 $Y=1.765
+ $X2=0 $Y2=0
cc_1101 N_A_2399_424#_c_1773_n N_VPWR_c_1813_n 0.0120466f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1102 N_A_2399_424#_M1011_g Q 0.00853833f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1103 N_A_2399_424#_M1011_g Q 0.00339956f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1104 N_A_2399_424#_c_1771_n Q 0.00791945f $X=12.93 $Y=1.765 $X2=0 $Y2=0
cc_1105 N_A_2399_424#_M1011_g Q 0.0228636f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1106 N_A_2399_424#_c_1793_p Q 0.0238691f $X=12.745 $Y=1.465 $X2=0 $Y2=0
cc_1107 N_A_2399_424#_c_1768_n N_VGND_c_2151_n 0.00917009f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1108 N_A_2399_424#_M1011_g N_VGND_c_2152_n 0.00647412f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1109 N_A_2399_424#_c_1767_n N_VGND_c_2152_n 0.00577732f $X=12.84 $Y=1.465
+ $X2=0 $Y2=0
cc_1110 N_A_2399_424#_c_1768_n N_VGND_c_2152_n 0.0504216f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1111 N_A_2399_424#_c_1793_p N_VGND_c_2152_n 0.0209147f $X=12.745 $Y=1.465
+ $X2=0 $Y2=0
cc_1112 N_A_2399_424#_c_1768_n N_VGND_c_2161_n 0.011066f $X=12.17 $Y=0.645 $X2=0
+ $Y2=0
cc_1113 N_A_2399_424#_M1011_g N_VGND_c_2162_n 0.00434272f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1114 N_A_2399_424#_M1011_g N_VGND_c_2163_n 0.00828941f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1115 N_A_2399_424#_c_1768_n N_VGND_c_2163_n 0.00915947f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1116 N_VPWR_c_1814_n N_A_300_464#_c_1982_n 0.0195202f $X=0.78 $Y=2.465 $X2=0
+ $Y2=0
cc_1117 N_VPWR_c_1830_n N_A_300_464#_c_1982_n 0.0471959f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1118 N_VPWR_c_1813_n N_A_300_464#_c_1982_n 0.0392475f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1119 N_VPWR_M1006_d N_A_300_464#_c_2001_n 0.0110267f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1120 N_VPWR_c_1815_n N_A_300_464#_c_2001_n 0.0214041f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1121 N_VPWR_c_1813_n N_A_300_464#_c_2001_n 0.0189567f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1122 N_VPWR_M1022_d N_A_300_464#_c_1984_n 0.0046335f $X=4.72 $Y=1.84 $X2=0
+ $Y2=0
cc_1123 N_VPWR_c_1816_n N_A_300_464#_c_1984_n 0.0166996f $X=4.87 $Y=2.815 $X2=0
+ $Y2=0
cc_1124 N_VPWR_c_1813_n N_A_300_464#_c_1984_n 0.0527404f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1125 N_VPWR_M1006_d N_A_300_464#_c_1985_n 8.56696e-19 $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1126 N_VPWR_c_1813_n N_A_300_464#_c_1985_n 0.00759345f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1127 N_VPWR_c_1831_n N_A_300_464#_c_1986_n 0.00535093f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_1128 N_VPWR_c_1813_n N_A_300_464#_c_1986_n 0.00675054f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1129 N_VPWR_c_1815_n N_A_300_464#_c_1990_n 0.00906624f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1130 N_VPWR_c_1815_n N_A_300_464#_c_1991_n 0.0176069f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1131 N_VPWR_c_1823_n N_A_300_464#_c_1991_n 0.0145459f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1132 N_VPWR_c_1813_n N_A_300_464#_c_1991_n 0.012028f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1133 N_VPWR_c_1822_n Q 0.0779559f $X=12.705 $Y=1.985 $X2=0 $Y2=0
cc_1134 N_VPWR_c_1833_n Q 0.0112891f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1135 N_VPWR_c_1813_n Q 0.00934413f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1136 N_A_300_464#_c_2001_n A_538_464# 0.00902149f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1137 N_A_300_464#_M1013_d N_noxref_24_c_2273_n 0.0106902f $X=1.95 $Y=0.405
+ $X2=0 $Y2=0
cc_1138 N_A_300_464#_c_1975_n N_noxref_24_c_2273_n 0.0460795f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1139 N_A_300_464#_c_1981_n N_noxref_24_c_2273_n 0.0239176f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1140 Q N_VGND_c_2152_n 0.0293763f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1141 Q N_VGND_c_2162_n 0.0145639f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1142 Q N_VGND_c_2163_n 0.0119984f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1143 N_VGND_c_2148_n N_noxref_24_c_2273_n 0.0231211f $X=3.87 $Y=0.565 $X2=0
+ $Y2=0
cc_1144 N_VGND_c_2153_n N_noxref_24_c_2273_n 0.142328f $X=3.785 $Y=0 $X2=0 $Y2=0
cc_1145 N_VGND_c_2163_n N_noxref_24_c_2273_n 0.0819703f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1146 N_VGND_c_2147_n N_noxref_24_c_2274_n 0.0259562f $X=0.71 $Y=0.65 $X2=0
+ $Y2=0
cc_1147 N_VGND_c_2153_n N_noxref_24_c_2274_n 0.0225398f $X=3.785 $Y=0 $X2=0
+ $Y2=0
cc_1148 N_VGND_c_2163_n N_noxref_24_c_2274_n 0.0125704f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1149 N_noxref_24_c_2273_n noxref_25 0.00198134f $X=3.09 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1150 N_noxref_24_c_2273_n noxref_26 0.00226367f $X=3.09 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
