* File: sky130_fd_sc_hs__fah_1.pex.spice
* Created: Thu Aug 27 20:46:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__FAH_1%CI 1 3 4 6 7 11
c40 11 0 1.05236e-19 $X=1.17 $Y=1.575
r41 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.575 $X2=1.17 $Y2=1.575
r42 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=1.665 $X2=1.17
+ $Y2=1.575
r43 4 10 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.185 $Y=1.825
+ $X2=1.17 $Y2=1.575
r44 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.185 $Y=1.825
+ $X2=1.185 $Y2=2.4
r45 1 10 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.08 $Y=1.41
+ $X2=1.17 $Y2=1.575
r46 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.08 $Y=1.41 $X2=1.08
+ $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_83_21# 1 2 10 11 12 13 15 16 17 19 25 30 31
+ 32 33 34 35 37 38 39 40 43 44 45 46 48 53 57 61 67
c189 53 0 1.16902e-20 $X=4.37 $Y=2.255
c190 46 0 2.4784e-20 $X=5.885 $Y=0.68
c191 34 0 3.05634e-20 $X=3.155 $Y=2.28
c192 31 0 3.93812e-19 $X=2.01 $Y=1.86
c193 25 0 1.37092e-19 $X=1.735 $Y=1.31
r194 61 64 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.05 $Y=0.68
+ $X2=6.05 $Y2=0.775
r195 57 59 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.96 $Y=0.68
+ $X2=4.96 $Y2=0.84
r196 53 55 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.37 $Y=2.255
+ $X2=4.37 $Y2=2.37
r197 48 50 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.24 $Y=2.28 $X2=3.24
+ $Y2=2.37
r198 47 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0.68
+ $X2=4.96 $Y2=0.68
r199 46 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.885 $Y=0.68
+ $X2=6.05 $Y2=0.68
r200 46 47 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.885 $Y=0.68
+ $X2=5.045 $Y2=0.68
r201 44 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=0.84
+ $X2=4.96 $Y2=0.84
r202 44 45 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.875 $Y=0.84
+ $X2=4.285 $Y2=0.84
r203 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=0.755
+ $X2=4.285 $Y2=0.84
r204 42 43 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.2 $Y=0.425
+ $X2=4.2 $Y2=0.755
r205 41 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.37
+ $X2=3.24 $Y2=2.37
r206 40 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=2.37
+ $X2=4.37 $Y2=2.37
r207 40 41 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=4.205 $Y=2.37
+ $X2=3.325 $Y2=2.37
r208 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.115 $Y=0.34
+ $X2=4.2 $Y2=0.425
r209 38 39 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.115 $Y=0.34
+ $X2=2.765 $Y2=0.34
r210 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.68 $Y=0.425
+ $X2=2.765 $Y2=0.34
r211 36 37 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.68 $Y=0.425
+ $X2=2.68 $Y2=0.9
r212 34 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=2.28
+ $X2=3.24 $Y2=2.28
r213 34 35 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=3.155 $Y=2.28
+ $X2=2.175 $Y2=2.28
r214 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.595 $Y=0.985
+ $X2=2.68 $Y2=0.9
r215 32 33 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.595 $Y=0.985
+ $X2=2.175 $Y2=0.985
r216 31 67 46.971 $w=5.15e-07 $l=1.65e-07 $layer=POLY_cond $X=1.917 $Y=1.86
+ $X2=1.917 $Y2=1.695
r217 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.01
+ $Y=1.86 $X2=2.01 $Y2=1.86
r218 28 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.01 $Y=2.195
+ $X2=2.175 $Y2=2.28
r219 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.01 $Y=2.195
+ $X2=2.01 $Y2=1.86
r220 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.01 $Y=1.07
+ $X2=2.175 $Y2=0.985
r221 27 30 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.01 $Y=1.07
+ $X2=2.01 $Y2=1.86
r222 23 25 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.62 $Y=1.31
+ $X2=1.735 $Y2=1.31
r223 20 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.735 $Y=1.385
+ $X2=1.735 $Y2=1.31
r224 20 67 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.735 $Y=1.385
+ $X2=1.735 $Y2=1.695
r225 19 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.62 $Y=1.235
+ $X2=1.62 $Y2=1.31
r226 18 19 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.62 $Y=0.255
+ $X2=1.62 $Y2=1.235
r227 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.545 $Y=0.18
+ $X2=1.62 $Y2=0.255
r228 16 17 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.545 $Y=0.18
+ $X2=0.565 $Y2=0.18
r229 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r230 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.675
+ $X2=0.505 $Y2=1.765
r231 11 22 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=1.375
r232 11 12 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=1.675
r233 10 22 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.49 $Y=0.93
+ $X2=0.49 $Y2=1.375
r234 7 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.49 $Y=0.255
+ $X2=0.565 $Y2=0.18
r235 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.49 $Y=0.255
+ $X2=0.49 $Y2=0.93
r236 2 53 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=4.22
+ $Y=2.12 $X2=4.37 $Y2=2.255
r237 1 64 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=5.84
+ $Y=0.625 $X2=6.05 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_410_58# 1 2 9 11 12 13 15 17 18 19 21 23 25
+ 27 29 34 35 38 39
c137 34 0 3.59827e-20 $X=4.88 $Y=1.26
c138 9 0 3.12094e-19 $X=2.125 $Y=0.79
r139 38 39 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=2.465
+ $X2=6.33 $Y2=2.465
r140 33 35 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=1.26
+ $X2=5.13 $Y2=1.26
r141 33 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=1.26
+ $X2=4.88 $Y2=1.26
r142 30 41 12.7214 $w=3.41e-07 $l=9e-08 $layer=POLY_cond $X=2.69 $Y=1.47
+ $X2=2.69 $Y2=1.38
r143 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.47 $X2=2.665 $Y2=1.47
r144 27 39 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.215 $Y=2.405
+ $X2=6.33 $Y2=2.405
r145 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.13 $Y=2.32
+ $X2=5.215 $Y2=2.405
r146 24 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=1.425
+ $X2=5.13 $Y2=1.26
r147 24 25 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=5.13 $Y=1.425
+ $X2=5.13 $Y2=2.32
r148 23 34 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=3.945 $Y=1.18 $X2=4.88
+ $Y2=1.18
r149 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.86 $Y=1.095
+ $X2=3.945 $Y2=1.18
r150 20 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.86 $Y=0.765
+ $X2=3.86 $Y2=1.095
r151 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.775 $Y=0.68
+ $X2=3.86 $Y2=0.765
r152 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.775 $Y=0.68
+ $X2=3.105 $Y2=0.68
r153 17 29 14.8322 $w=2.92e-07 $l=4.42674e-07 $layer=LI1_cond $X=3.02 $Y=1.24
+ $X2=2.665 $Y2=1.437
r154 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=0.765
+ $X2=3.105 $Y2=0.68
r155 16 17 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.02 $Y=0.765
+ $X2=3.02 $Y2=1.24
r156 13 30 57.0643 $w=3.41e-07 $l=3.41358e-07 $layer=POLY_cond $X=2.79 $Y=1.765
+ $X2=2.69 $Y2=1.47
r157 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.79 $Y=1.765
+ $X2=2.79 $Y2=2.4
r158 11 41 22.0049 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.5 $Y=1.38
+ $X2=2.69 $Y2=1.38
r159 11 12 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.5 $Y=1.38 $X2=2.2
+ $Y2=1.38
r160 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=1.305
+ $X2=2.2 $Y2=1.38
r161 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.125 $Y=1.305
+ $X2=2.125 $Y2=0.79
r162 2 38 600 $w=1.7e-07 $l=6.80882e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=1.865 $X2=6.495 $Y2=2.475
r163 1 33 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=4.905
+ $Y=0.835 $X2=5.045 $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_231_132# 1 2 3 4 13 15 16 18 21 26 29 30 31
+ 33 37 40 41 43 46 47 49 50 52 54 55 56 60 65 66 68 69 71 77
c244 66 0 1.16902e-20 $X=4.175 $Y=1.52
c245 65 0 7.86143e-20 $X=4.175 $Y=1.52
c246 55 0 1.55643e-19 $X=1.5 $Y=1.95
c247 31 0 3.05363e-20 $X=3.46 $Y=2.71
c248 21 0 2.93543e-19 $X=1.505 $Y=1.155
r249 76 77 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.96 $Y=2.902
+ $X2=6.125 $Y2=2.902
r250 71 73 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.55 $Y=1.03 $X2=5.55
+ $Y2=1.12
r251 65 68 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.175 $Y=1.6
+ $X2=4.34 $Y2=1.6
r252 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.175
+ $Y=1.52 $X2=4.175 $Y2=1.52
r253 60 62 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.545 $Y=2.71
+ $X2=3.545 $Y2=2.99
r254 56 58 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.9 $Y=2.62 $X2=2.9
+ $Y2=2.71
r255 54 55 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.5 $Y=2.115
+ $X2=1.5 $Y2=1.95
r256 51 52 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.915 $Y=2.12
+ $X2=6.915 $Y2=2.905
r257 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.83 $Y=2.035
+ $X2=6.915 $Y2=2.12
r258 49 50 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.83 $Y=2.035
+ $X2=6.225 $Y2=2.035
r259 47 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.83 $Y=2.99
+ $X2=6.915 $Y2=2.905
r260 47 77 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.83 $Y=2.99
+ $X2=6.125 $Y2=2.99
r261 46 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.14 $Y=1.95
+ $X2=6.225 $Y2=2.035
r262 45 46 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=6.14 $Y=1.205
+ $X2=6.14 $Y2=1.95
r263 44 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=1.12
+ $X2=5.55 $Y2=1.12
r264 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.055 $Y=1.12
+ $X2=6.14 $Y2=1.205
r265 43 44 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.055 $Y=1.12
+ $X2=5.715 $Y2=1.12
r266 42 69 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=2.902
+ $X2=4.79 $Y2=2.902
r267 41 76 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=5.953 $Y=2.902
+ $X2=5.96 $Y2=2.902
r268 41 42 36.0097 $w=3.43e-07 $l=1.078e-06 $layer=LI1_cond $X=5.953 $Y=2.902
+ $X2=4.875 $Y2=2.902
r269 40 69 2.87242 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.79 $Y=2.73
+ $X2=4.79 $Y2=2.902
r270 39 40 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=4.79 $Y=1.765
+ $X2=4.79 $Y2=2.73
r271 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.705 $Y=1.68
+ $X2=4.79 $Y2=1.765
r272 37 68 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.705 $Y=1.68
+ $X2=4.34 $Y2=1.68
r273 34 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=2.99
+ $X2=3.545 $Y2=2.99
r274 33 69 3.6114 $w=2.57e-07 $l=1.23386e-07 $layer=LI1_cond $X=4.705 $Y=2.99
+ $X2=4.79 $Y2=2.902
r275 33 34 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=4.705 $Y=2.99
+ $X2=3.63 $Y2=2.99
r276 32 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=2.71
+ $X2=2.9 $Y2=2.71
r277 31 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=2.71
+ $X2=3.545 $Y2=2.71
r278 31 32 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.46 $Y=2.71
+ $X2=2.985 $Y2=2.71
r279 29 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=2.62
+ $X2=2.9 $Y2=2.62
r280 29 30 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.815 $Y=2.62
+ $X2=1.675 $Y2=2.62
r281 27 55 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.59 $Y=1.24
+ $X2=1.59 $Y2=1.95
r282 26 30 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=1.5 $Y=2.535
+ $X2=1.675 $Y2=2.62
r283 25 54 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=1.5 $Y=2.125 $X2=1.5
+ $Y2=2.115
r284 25 26 13.5 $w=3.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.5 $Y=2.125 $X2=1.5
+ $Y2=2.535
r285 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=1.155
+ $X2=1.59 $Y2=1.24
r286 21 23 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.505 $Y=1.155
+ $X2=1.31 $Y2=1.155
r287 20 66 81.236 $w=4.45e-07 $l=6.5e-07 $layer=POLY_cond $X=3.525 $Y=1.462
+ $X2=4.175 $Y2=1.462
r288 16 20 74.3954 $w=2.52e-07 $l=3.90415e-07 $layer=POLY_cond $X=3.435 $Y=1.81
+ $X2=3.345 $Y2=1.462
r289 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.435 $Y=1.81
+ $X2=3.435 $Y2=2.385
r290 13 20 50.2954 $w=2.52e-07 $l=3.06078e-07 $layer=POLY_cond $X=3.145 $Y=1.24
+ $X2=3.345 $Y2=1.462
r291 13 15 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.145 $Y=1.24
+ $X2=3.145 $Y2=0.84
r292 4 76 300 $w=1.7e-07 $l=9.77561e-07 $layer=licon1_PDIFF $count=2 $X=5.28
+ $Y=2.12 $X2=5.96 $Y2=2.815
r293 3 54 300 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=2 $X=1.26
+ $Y=1.9 $X2=1.41 $Y2=2.115
r294 2 71 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=5.41
+ $Y=0.625 $X2=5.55 $Y2=1.03
r295 1 23 182 $w=1.7e-07 $l=5.6723e-07 $layer=licon1_NDIFF $count=1 $X=1.155
+ $Y=0.66 $X2=1.31 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_811_379# 1 2 7 9 10 11 13 17 18 19 23 24 26
+ 28 31 33 34 36 41 42 46 49 50 53 56 57
c205 41 0 4.59067e-20 $X=5.785 $Y=1.54
r206 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.925 $Y=2.035
+ $X2=8.925 $Y2=2.035
r207 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r208 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r209 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.78 $Y=2.035
+ $X2=8.925 $Y2=2.035
r210 49 50 3.85519 $w=1.4e-07 $l=3.115e-06 $layer=MET1_cond $X=8.78 $Y=2.035
+ $X2=5.665 $Y2=2.035
r211 46 48 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=10.65 $Y=0.82
+ $X2=10.65 $Y2=1.05
r212 44 57 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=8.945 $Y=2.565
+ $X2=8.945 $Y2=2.035
r213 42 61 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.785 $Y=1.54
+ $X2=5.785 $Y2=1.715
r214 42 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.785 $Y=1.54
+ $X2=5.785 $Y2=1.375
r215 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.785
+ $Y=1.54 $X2=5.785 $Y2=1.54
r216 38 53 16.5351 $w=2.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.52 $Y=1.705
+ $X2=5.52 $Y2=2.035
r217 37 41 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=5.52 $Y=1.54
+ $X2=5.785 $Y2=1.54
r218 37 38 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.52 $Y=1.54
+ $X2=5.52 $Y2=1.705
r219 36 48 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=10.73 $Y=2.565
+ $X2=10.73 $Y2=1.05
r220 34 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.11 $Y=2.65
+ $X2=8.945 $Y2=2.565
r221 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.645 $Y=2.65
+ $X2=10.73 $Y2=2.565
r222 33 34 100.144 $w=1.68e-07 $l=1.535e-06 $layer=LI1_cond $X=10.645 $Y=2.65
+ $X2=9.11 $Y2=2.65
r223 29 31 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.655 $Y=1.625
+ $X2=4.83 $Y2=1.625
r224 26 28 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.27 $Y=1.79
+ $X2=6.27 $Y2=2.285
r225 25 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.715
+ $X2=5.785 $Y2=1.715
r226 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.195 $Y=1.715
+ $X2=6.27 $Y2=1.79
r227 24 25 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=6.195 $Y=1.715
+ $X2=5.95 $Y2=1.715
r228 23 60 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.765 $Y=0.945
+ $X2=5.765 $Y2=1.375
r229 20 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.765 $Y=0.255
+ $X2=5.765 $Y2=0.945
r230 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.69 $Y=0.18
+ $X2=5.765 $Y2=0.255
r231 18 19 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.69 $Y=0.18
+ $X2=4.905 $Y2=0.18
r232 15 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.83 $Y=1.55
+ $X2=4.83 $Y2=1.625
r233 15 17 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.83 $Y=1.55
+ $X2=4.83 $Y2=1.155
r234 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.83 $Y=0.255
+ $X2=4.905 $Y2=0.18
r235 14 17 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=4.83 $Y=0.255
+ $X2=4.83 $Y2=1.155
r236 12 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.655 $Y=1.7
+ $X2=4.655 $Y2=1.625
r237 12 13 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.655 $Y=1.7
+ $X2=4.655 $Y2=1.895
r238 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.58 $Y=1.97
+ $X2=4.655 $Y2=1.895
r239 10 11 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.58 $Y=1.97
+ $X2=4.22 $Y2=1.97
r240 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.145 $Y=2.045
+ $X2=4.22 $Y2=1.97
r241 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.145 $Y=2.045
+ $X2=4.145 $Y2=2.54
r242 2 57 300 $w=1.7e-07 $l=2.88141e-07 $layer=licon1_PDIFF $count=2 $X=8.745
+ $Y=1.87 $X2=8.945 $Y2=2.075
r243 1 46 182 $w=1.7e-07 $l=6.20806e-07 $layer=licon1_NDIFF $count=1 $X=10.18
+ $Y=0.47 $X2=10.65 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_1023_379# 1 2 10 13 15 16 17 19 20 21 23 24
+ 25 26 29 32 35 38 39 43 47 53 55 56 57 58 61 64 65 70 73
c215 65 0 3.01025e-19 $X=11.1 $Y=1.665
c216 61 0 1.03145e-19 $X=6.96 $Y=1.665
c217 38 0 1.45758e-19 $X=6.9 $Y=0.875
c218 21 0 2.11227e-20 $X=6.34 $Y=1.325
r219 65 74 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.1 $Y=1.665
+ $X2=11.1 $Y2=1.78
r220 65 73 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.1 $Y=1.665
+ $X2=11.1 $Y2=1.55
r221 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.1 $Y=1.665
+ $X2=11.1 $Y2=1.665
r222 61 70 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.55
r223 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.665
r224 58 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=1.665
+ $X2=6.96 $Y2=1.665
r225 57 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.955 $Y=1.665
+ $X2=11.1 $Y2=1.665
r226 57 58 4.76484 $w=1.4e-07 $l=3.85e-06 $layer=MET1_cond $X=10.955 $Y=1.665
+ $X2=7.105 $Y2=1.665
r227 55 70 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=6.955 $Y=1.38
+ $X2=6.955 $Y2=1.55
r228 53 74 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=11.07 $Y=1.98
+ $X2=11.07 $Y2=1.78
r229 49 73 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=11.07 $Y=0.425
+ $X2=11.07 $Y2=1.55
r230 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.985 $Y=0.34
+ $X2=11.07 $Y2=0.425
r231 47 56 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=10.985 $Y=0.34
+ $X2=9.385 $Y2=0.34
r232 43 56 5.72867 $w=1.93e-07 $l=9.7e-08 $layer=LI1_cond $X=9.288 $Y=0.352
+ $X2=9.385 $Y2=0.352
r233 43 45 8.41772 $w=1.93e-07 $l=1.48e-07 $layer=LI1_cond $X=9.288 $Y=0.352
+ $X2=9.14 $Y2=0.352
r234 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.9
+ $Y=0.875 $X2=6.9 $Y2=0.875
r235 36 55 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.9 $Y=1.215
+ $X2=6.9 $Y2=1.38
r236 36 38 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.9 $Y=1.215
+ $X2=6.9 $Y2=0.875
r237 34 39 61.826 $w=3.5e-07 $l=3.75e-07 $layer=POLY_cond $X=6.91 $Y=1.25
+ $X2=6.91 $Y2=0.875
r238 34 35 12.4285 $w=2.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.91 $Y=1.25
+ $X2=6.925 $Y2=1.325
r239 30 32 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=5.205 $Y=1.97
+ $X2=5.335 $Y2=1.97
r240 27 29 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.025 $Y=2.78
+ $X2=7.025 $Y2=2.285
r241 26 29 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.025 $Y=1.79
+ $X2=7.025 $Y2=2.285
r242 24 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.025 $Y=2.87
+ $X2=7.025 $Y2=2.78
r243 24 25 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=7.025 $Y=2.87
+ $X2=7.025 $Y2=3.075
r244 23 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.025 $Y=1.7
+ $X2=7.025 $Y2=1.79
r245 22 35 12.4285 $w=2.65e-07 $l=1.32288e-07 $layer=POLY_cond $X=7.025 $Y=1.4
+ $X2=6.925 $Y2=1.325
r246 22 23 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=7.025 $Y=1.4
+ $X2=7.025 $Y2=1.7
r247 20 35 13.6393 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.735 $Y=1.325
+ $X2=6.925 $Y2=1.325
r248 20 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.735 $Y=1.325
+ $X2=6.34 $Y2=1.325
r249 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.265 $Y=1.25
+ $X2=6.34 $Y2=1.325
r250 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.265 $Y=1.25
+ $X2=6.265 $Y2=0.855
r251 15 25 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.935 $Y=3.15
+ $X2=7.025 $Y2=3.075
r252 15 16 840.936 $w=1.5e-07 $l=1.64e-06 $layer=POLY_cond $X=6.935 $Y=3.15
+ $X2=5.295 $Y2=3.15
r253 11 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.335 $Y=1.895
+ $X2=5.335 $Y2=1.97
r254 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.335 $Y=1.895
+ $X2=5.335 $Y2=0.945
r255 8 16 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=5.205 $Y=3.035
+ $X2=5.295 $Y2=3.15
r256 8 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.205 $Y=3.035
+ $X2=5.205 $Y2=2.54
r257 7 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.205 $Y=2.045
+ $X2=5.205 $Y2=1.97
r258 7 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.205 $Y=2.045
+ $X2=5.205 $Y2=2.54
r259 2 53 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=10.92
+ $Y=1.84 $X2=11.07 $Y2=1.98
r260 1 45 182 $w=1.7e-07 $l=3.48569e-07 $layer=licon1_NDIFF $count=1 $X=8.84
+ $Y=0.47 $X2=9.14 $Y2=0.365
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_879_55# 1 2 3 10 12 15 17 19 20 22 24 25 27
+ 31 36 38 41 44 45 49 55 56 57 58 63 65 67 69 75
c194 27 0 3.59827e-20 $X=7.235 $Y=0.34
c195 10 0 1.50564e-19 $X=8.67 $Y=1.795
r196 68 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.31 $Y=1.385
+ $X2=10.475 $Y2=1.385
r197 68 72 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=10.31 $Y=1.385
+ $X2=10.105 $Y2=1.385
r198 67 69 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.31 $Y=1.385
+ $X2=10.31 $Y2=1.22
r199 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.31
+ $Y=1.385 $X2=10.31 $Y2=1.385
r200 60 63 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=8.675 $Y=1.545
+ $X2=8.89 $Y2=1.545
r201 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.675
+ $Y=1.545 $X2=8.675 $Y2=1.545
r202 56 58 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=7.415 $Y=1.95
+ $X2=7.415 $Y2=1.13
r203 55 56 6.19221 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=7.335 $Y=2.05
+ $X2=7.335 $Y2=1.95
r204 49 52 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.58 $Y=0.34 $X2=4.58
+ $Y2=0.42
r205 47 69 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.23 $Y=0.79
+ $X2=10.23 $Y2=1.22
r206 46 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.975 $Y=0.705
+ $X2=8.89 $Y2=0.705
r207 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.145 $Y=0.705
+ $X2=10.23 $Y2=0.79
r208 45 46 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=10.145 $Y=0.705
+ $X2=8.975 $Y2=0.705
r209 44 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.89 $Y=1.38
+ $X2=8.89 $Y2=1.545
r210 43 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.89 $Y=0.79
+ $X2=8.89 $Y2=0.705
r211 43 44 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.89 $Y=0.79
+ $X2=8.89 $Y2=1.38
r212 42 57 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.565 $Y=0.705
+ $X2=7.4 $Y2=0.705
r213 41 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.805 $Y=0.705
+ $X2=8.89 $Y2=0.705
r214 41 42 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=8.805 $Y=0.705
+ $X2=7.565 $Y2=0.705
r215 38 58 7.25185 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.4 $Y=0.965
+ $X2=7.4 $Y2=1.13
r216 37 57 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=0.79 $X2=7.4
+ $Y2=0.705
r217 37 38 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.4 $Y=0.79
+ $X2=7.4 $Y2=0.965
r218 34 57 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=0.62 $X2=7.4
+ $Y2=0.705
r219 34 36 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.4 $Y=0.62
+ $X2=7.4 $Y2=0.515
r220 33 36 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.4 $Y=0.425 $X2=7.4
+ $Y2=0.515
r221 29 55 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=7.335 $Y=2.115
+ $X2=7.335 $Y2=2.05
r222 29 31 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=7.335 $Y=2.115
+ $X2=7.335 $Y2=2.76
r223 28 49 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.705 $Y=0.34
+ $X2=4.58 $Y2=0.34
r224 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.235 $Y=0.34
+ $X2=7.4 $Y2=0.425
r225 27 28 165.059 $w=1.68e-07 $l=2.53e-06 $layer=LI1_cond $X=7.235 $Y=0.34
+ $X2=4.705 $Y2=0.34
r226 22 25 114.876 $w=1.8e-07 $l=2.9e-07 $layer=POLY_cond $X=10.845 $Y=1.765
+ $X2=10.845 $Y2=1.475
r227 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.845 $Y=1.765
+ $X2=10.845 $Y2=2.26
r228 20 25 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.755 $Y=1.475
+ $X2=10.845 $Y2=1.475
r229 20 75 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.755 $Y=1.475
+ $X2=10.475 $Y2=1.475
r230 17 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.105 $Y=1.22
+ $X2=10.105 $Y2=1.385
r231 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.105 $Y=1.22
+ $X2=10.105 $Y2=0.79
r232 13 61 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=8.765 $Y=1.38
+ $X2=8.675 $Y2=1.545
r233 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.765 $Y=1.38
+ $X2=8.765 $Y2=0.79
r234 10 61 52.2586 $w=2.99e-07 $l=2.52488e-07 $layer=POLY_cond $X=8.67 $Y=1.795
+ $X2=8.675 $Y2=1.545
r235 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.67 $Y=1.795
+ $X2=8.67 $Y2=2.29
r236 3 55 300 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_PDIFF $count=2 $X=7.1
+ $Y=1.865 $X2=7.335 $Y2=2.05
r237 3 31 600 $w=1.7e-07 $l=1.00566e-06 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.865 $X2=7.335 $Y2=2.76
r238 2 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.255
+ $Y=0.37 $X2=7.4 $Y2=0.515
r239 1 52 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.395
+ $Y=0.275 $X2=4.54 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%B 1 3 6 8 11 12 13 15 16 17 18 21 22 24 26 29
+ 32 33 34 35 38 39 40 42 43 50
c157 43 0 1.50564e-19 $X=9.36 $Y=1.295
c158 38 0 1.04105e-19 $X=11.295 $Y=2.26
c159 8 0 1.01602e-19 $X=8.055 $Y=1.635
c160 6 0 1.45758e-19 $X=7.615 $Y=0.74
c161 1 0 1.03145e-19 $X=7.56 $Y=1.71
r162 48 50 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=9.31 $Y=1.385
+ $X2=9.515 $Y2=1.385
r163 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.31
+ $Y=1.385 $X2=9.31 $Y2=1.385
r164 45 48 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=9.17 $Y=1.385
+ $X2=9.31 $Y2=1.385
r165 43 49 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.31 $Y=1.295
+ $X2=9.31 $Y2=1.385
r166 41 42 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=11.292 $Y=1.35
+ $X2=11.292 $Y2=1.5
r167 36 38 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=11.295 $Y=2.76
+ $X2=11.295 $Y2=2.26
r168 35 38 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.295 $Y=1.765
+ $X2=11.295 $Y2=2.26
r169 33 36 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.295 $Y=2.85
+ $X2=11.295 $Y2=2.76
r170 33 34 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=11.295 $Y=2.85
+ $X2=11.295 $Y2=3.075
r171 32 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.295 $Y=1.675
+ $X2=11.295 $Y2=1.765
r172 32 42 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=11.295 $Y=1.675
+ $X2=11.295 $Y2=1.5
r173 29 41 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.275 $Y=0.79
+ $X2=11.275 $Y2=1.35
r174 24 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.515 $Y=1.22
+ $X2=9.515 $Y2=1.385
r175 24 26 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.515 $Y=1.22
+ $X2=9.515 $Y2=0.79
r176 23 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.26 $Y=3.15 $X2=9.17
+ $Y2=3.15
r177 22 34 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=11.205 $Y=3.15
+ $X2=11.295 $Y2=3.075
r178 22 23 997.33 $w=1.5e-07 $l=1.945e-06 $layer=POLY_cond $X=11.205 $Y=3.15
+ $X2=9.26 $Y2=3.15
r179 19 21 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.17 $Y=2.785
+ $X2=9.17 $Y2=2.29
r180 18 21 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.17 $Y=1.795
+ $X2=9.17 $Y2=2.29
r181 17 40 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.17 $Y=3.075
+ $X2=9.17 $Y2=3.15
r182 16 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.17 $Y=2.875
+ $X2=9.17 $Y2=2.785
r183 16 17 77.7419 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=9.17 $Y=2.875
+ $X2=9.17 $Y2=3.075
r184 15 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.17 $Y=1.705
+ $X2=9.17 $Y2=1.795
r185 14 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.17 $Y=1.55
+ $X2=9.17 $Y2=1.385
r186 14 15 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=9.17 $Y=1.55
+ $X2=9.17 $Y2=1.705
r187 12 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.08 $Y=3.15 $X2=9.17
+ $Y2=3.15
r188 12 13 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=9.08 $Y=3.15
+ $X2=8.205 $Y2=3.15
r189 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.13 $Y=3.075
+ $X2=8.205 $Y2=3.15
r190 10 11 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=8.13 $Y=1.71
+ $X2=8.13 $Y2=3.075
r191 9 39 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=7.69 $Y=1.635
+ $X2=7.58 $Y2=1.635
r192 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.055 $Y=1.635
+ $X2=8.13 $Y2=1.71
r193 8 9 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=8.055 $Y=1.635
+ $X2=7.69 $Y2=1.635
r194 4 39 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=7.615 $Y=1.56
+ $X2=7.58 $Y2=1.635
r195 4 6 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.615 $Y=1.56
+ $X2=7.615 $Y2=0.74
r196 1 39 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=7.56 $Y=1.71
+ $X2=7.58 $Y2=1.635
r197 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.56 $Y=1.71
+ $X2=7.56 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_2342_48# 1 2 9 10 12 14 15 16 20 24 28 32 35
+ 36 37
c81 28 0 1.0013e-19 $X=12.415 $Y=1.215
c82 14 0 1.96919e-19 $X=11.89 $Y=1.385
r83 35 36 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=13.65 $Y=2.135
+ $X2=13.65 $Y2=1.97
r84 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.415
+ $Y=1.385 $X2=12.415 $Y2=1.385
r85 28 31 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=12.415 $Y=1.215
+ $X2=12.415 $Y2=1.385
r86 26 37 3.55013 $w=2.62e-07 $l=1.28662e-07 $layer=LI1_cond $X=13.745 $Y=1.3
+ $X2=13.652 $Y2=1.215
r87 26 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.745 $Y=1.3
+ $X2=13.745 $Y2=1.97
r88 22 37 3.55013 $w=2.62e-07 $l=8.5e-08 $layer=LI1_cond $X=13.652 $Y=1.13
+ $X2=13.652 $Y2=1.215
r89 22 24 19.9649 $w=3.53e-07 $l=6.15e-07 $layer=LI1_cond $X=13.652 $Y=1.13
+ $X2=13.652 $Y2=0.515
r90 18 35 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=13.65 $Y=2.15
+ $X2=13.65 $Y2=2.135
r91 18 20 21.2882 $w=3.58e-07 $l=6.65e-07 $layer=LI1_cond $X=13.65 $Y=2.15
+ $X2=13.65 $Y2=2.815
r92 17 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.58 $Y=1.215
+ $X2=12.415 $Y2=1.215
r93 16 37 2.9446 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=13.475 $Y=1.215
+ $X2=13.652 $Y2=1.215
r94 16 17 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=13.475 $Y=1.215
+ $X2=12.58 $Y2=1.215
r95 14 32 91.8022 $w=3.3e-07 $l=5.25e-07 $layer=POLY_cond $X=11.89 $Y=1.385
+ $X2=12.415 $Y2=1.385
r96 14 15 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.8 $Y=1.385
+ $X2=11.8 $Y2=1.22
r97 10 14 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=11.8 $Y=1.765
+ $X2=11.8 $Y2=1.385
r98 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.8 $Y=1.765
+ $X2=11.8 $Y2=2.4
r99 9 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.785 $Y=0.74
+ $X2=11.785 $Y2=1.22
r100 2 35 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=13.485
+ $Y=1.96 $X2=13.635 $Y2=2.135
r101 2 20 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=13.485
+ $Y=1.96 $X2=13.635 $Y2=2.815
r102 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.5
+ $Y=0.37 $X2=13.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A 3 5 7 8 10 13 15 21 22
c48 22 0 1.0013e-19 $X=13.41 $Y=1.677
r49 22 23 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=13.41 $Y=1.677
+ $X2=13.425 $Y2=1.677
r50 20 22 10.9253 $w=3.75e-07 $l=8.5e-08 $layer=POLY_cond $X=13.325 $Y=1.677
+ $X2=13.41 $Y2=1.677
r51 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.325
+ $Y=1.635 $X2=13.325 $Y2=1.635
r52 18 20 53.3413 $w=3.75e-07 $l=4.15e-07 $layer=POLY_cond $X=12.91 $Y=1.677
+ $X2=13.325 $Y2=1.677
r53 17 18 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=12.895 $Y=1.677
+ $X2=12.91 $Y2=1.677
r54 15 21 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=13.2 $Y=1.635
+ $X2=13.325 $Y2=1.635
r55 11 23 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.425 $Y=1.47
+ $X2=13.425 $Y2=1.677
r56 11 13 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=13.425 $Y=1.47
+ $X2=13.425 $Y2=0.69
r57 8 22 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=13.41 $Y=1.885
+ $X2=13.41 $Y2=1.677
r58 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=13.41 $Y=1.885
+ $X2=13.41 $Y2=2.46
r59 5 18 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=12.91 $Y=1.885
+ $X2=12.91 $Y2=1.677
r60 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.91 $Y=1.885
+ $X2=12.91 $Y2=2.46
r61 1 17 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.895 $Y=1.47
+ $X2=12.895 $Y2=1.677
r62 1 3 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=12.895 $Y=1.47
+ $X2=12.895 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%SUM 1 2 7 8 9 10 11 18
r18 10 11 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=2.405
+ $X2=0.277 $Y2=2.775
r19 9 10 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=0.277 $Y=1.985
+ $X2=0.277 $Y2=2.405
r20 8 9 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.985
r21 7 8 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.665
r22 7 18 20.2968 $w=3.33e-07 $l=5.9e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=0.705
r23 2 11 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r24 2 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r25 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.56 $X2=0.275 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%VPWR 1 2 3 4 5 20 24 28 31 36 43 44 45 47 55
+ 67 73 74 77 80 87 90
c132 80 0 3.05634e-20 $X=3.11 $Y=3.05
r133 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r134 87 88 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r135 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r136 74 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r137 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r138 71 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.3 $Y=3.33
+ $X2=13.175 $Y2=3.33
r139 71 73 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=13.3 $Y=3.33
+ $X2=13.68 $Y2=3.33
r140 70 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r141 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r142 67 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.05 $Y=3.33
+ $X2=13.175 $Y2=3.33
r143 67 69 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=13.05 $Y=3.33
+ $X2=12.72 $Y2=3.33
r144 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r145 66 88 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=7.92 $Y2=3.33
r146 65 66 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r147 63 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8 $Y=3.33 $X2=7.835
+ $Y2=3.33
r148 63 65 245.305 $w=1.68e-07 $l=3.76e-06 $layer=LI1_cond $X=8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r149 62 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r150 61 62 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r151 59 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r152 58 61 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r153 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r154 56 58 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.29 $Y=3.33
+ $X2=3.6 $Y2=3.33
r155 55 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.67 $Y=3.33
+ $X2=7.835 $Y2=3.33
r156 55 61 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.67 $Y=3.33
+ $X2=7.44 $Y2=3.33
r157 54 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r158 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r159 51 54 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r160 51 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r161 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r162 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r163 48 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r164 48 50 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r165 47 56 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=3.112 $Y=3.33
+ $X2=3.29 $Y2=3.33
r166 47 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r167 47 80 9.08969 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=3.112 $Y=3.33
+ $X2=3.112 $Y2=3.05
r168 47 53 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=3.33
+ $X2=2.64 $Y2=3.33
r169 45 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r170 45 59 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=3.6 $Y2=3.33
r171 43 65 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.95 $Y=3.33
+ $X2=11.76 $Y2=3.33
r172 43 44 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.95 $Y=3.33
+ $X2=12.12 $Y2=3.33
r173 42 69 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=12.29 $Y=3.33
+ $X2=12.72 $Y2=3.33
r174 42 44 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.29 $Y=3.33
+ $X2=12.12 $Y2=3.33
r175 36 39 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=13.175 $Y=2.135
+ $X2=13.175 $Y2=2.815
r176 34 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.175 $Y=3.245
+ $X2=13.175 $Y2=3.33
r177 34 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=13.175 $Y=3.245
+ $X2=13.175 $Y2=2.815
r178 31 33 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=12.12 $Y=2.615
+ $X2=12.12 $Y2=2.955
r179 29 44 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=12.12 $Y=3.245
+ $X2=12.12 $Y2=3.33
r180 29 33 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=12.12 $Y=3.245
+ $X2=12.12 $Y2=2.955
r181 28 41 8.27282 $w=3.4e-07 $l=2.25e-07 $layer=LI1_cond $X=12.12 $Y=2.5
+ $X2=12.12 $Y2=2.275
r182 28 31 3.89797 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=12.12 $Y=2.5
+ $X2=12.12 $Y2=2.615
r183 24 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.835 $Y=1.93
+ $X2=7.835 $Y2=2.76
r184 22 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.835 $Y=3.245
+ $X2=7.835 $Y2=3.33
r185 22 27 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=7.835 $Y=3.245
+ $X2=7.835 $Y2=2.76
r186 18 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r187 18 20 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r188 5 39 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=12.985
+ $Y=1.96 $X2=13.135 $Y2=2.815
r189 5 36 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=12.985
+ $Y=1.96 $X2=13.135 $Y2=2.135
r190 4 41 600 $w=1.7e-07 $l=5.41872e-07 $layer=licon1_PDIFF $count=1 $X=11.875
+ $Y=1.84 $X2=12.115 $Y2=2.275
r191 4 33 600 $w=1.7e-07 $l=1.22916e-06 $layer=licon1_PDIFF $count=1 $X=11.875
+ $Y=1.84 $X2=12.115 $Y2=2.955
r192 4 31 600 $w=1.7e-07 $l=8.86919e-07 $layer=licon1_PDIFF $count=1 $X=11.875
+ $Y=1.84 $X2=12.115 $Y2=2.615
r193 3 27 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.785 $X2=7.835 $Y2=2.76
r194 3 24 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.785 $X2=7.835 $Y2=1.93
r195 2 80 600 $w=1.7e-07 $l=1.32686e-06 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=1.84 $X2=3.11 $Y2=3.05
r196 1 20 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%COUT 1 2 8 9 10 12 14 17 20 21 23
c75 17 0 1.15685e-19 $X=1.07 $Y=2.035
c76 12 0 1.72891e-19 $X=1.07 $Y=2.905
r77 23 28 7.38421 $w=3.8e-07 $l=2.3e-07 $layer=LI1_cond $X=1.68 $Y=0.65 $X2=1.91
+ $Y2=0.65
r78 20 21 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=2.975
+ $X2=2.315 $Y2=2.975
r79 15 17 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.75 $Y=2.035
+ $X2=1.07 $Y2=2.035
r80 14 21 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=1.155 $Y=2.99
+ $X2=2.315 $Y2=2.99
r81 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=2.905
+ $X2=1.155 $Y2=2.99
r82 11 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=2.12
+ $X2=1.07 $Y2=2.035
r83 11 12 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.07 $Y=2.12
+ $X2=1.07 $Y2=2.905
r84 9 23 9.3947 $w=3.8e-07 $l=2.43926e-07 $layer=LI1_cond $X=1.505 $Y=0.815
+ $X2=1.68 $Y2=0.65
r85 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.505 $Y=0.815
+ $X2=0.835 $Y2=0.815
r86 8 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.95 $X2=0.75
+ $Y2=2.035
r87 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.75 $Y=0.9
+ $X2=0.835 $Y2=0.815
r88 7 8 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=0.75 $Y=0.9 $X2=0.75
+ $Y2=1.95
r89 2 20 600 $w=1.7e-07 $l=1.19029e-06 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.84 $X2=2.48 $Y2=2.96
r90 1 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.42 $X2=1.91 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_644_104# 1 2 3 11 14 17 20 21 27 28 31
c98 31 0 3.05363e-20 $X=3.36 $Y=1.855
c99 21 0 7.86143e-20 $X=3.265 $Y=1.665
r100 31 33 13.9377 $w=3.37e-07 $l=3.85e-07 $layer=LI1_cond $X=3.36 $Y=1.855
+ $X2=3.745 $Y2=1.855
r101 28 35 6.65862 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=6.495 $Y=1.665
+ $X2=6.495 $Y2=1.55
r102 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r103 24 31 8.68843 $w=3.37e-07 $l=2.4e-07 $layer=LI1_cond $X=3.12 $Y=1.855
+ $X2=3.36 $Y2=1.855
r104 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r105 21 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r106 20 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=6.48 $Y2=1.665
r107 20 21 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=3.265 $Y2=1.665
r108 17 19 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=1.02
+ $X2=3.44 $Y2=1.185
r109 14 35 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.48 $Y=0.875
+ $X2=6.48 $Y2=1.55
r110 11 31 4.74843 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.36 $Y=1.58
+ $X2=3.36 $Y2=1.855
r111 11 19 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.36 $Y=1.58
+ $X2=3.36 $Y2=1.185
r112 3 33 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.51
+ $Y=1.885 $X2=3.745 $Y2=2.03
r113 2 14 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.535 $X2=6.48 $Y2=0.875
r114 1 17 182 $w=1.7e-07 $l=6e-07 $layer=licon1_NDIFF $count=1 $X=3.22 $Y=0.52
+ $X2=3.44 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_1660_374# 1 2 3 4 16 17 18 19 22 25 32 35 36
c91 32 0 1.01602e-19 $X=8.47 $Y=1.045
r92 35 36 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=8.39 $Y=2.045
+ $X2=8.39 $Y2=1.88
r93 29 32 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=8.255 $Y=1.085
+ $X2=8.47 $Y2=1.085
r94 28 37 5.67621 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=11.572 $Y=0.965
+ $X2=11.572 $Y2=1.13
r95 25 28 15.4806 $w=3.33e-07 $l=4.5e-07 $layer=LI1_cond $X=11.572 $Y=0.515
+ $X2=11.572 $Y2=0.965
r96 20 22 29.7038 $w=3.53e-07 $l=9.15e-07 $layer=LI1_cond $X=11.562 $Y=2.905
+ $X2=11.562 $Y2=1.99
r97 19 37 5.79584 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=11.562 $Y=1.307
+ $X2=11.562 $Y2=1.13
r98 19 22 22.1724 $w=3.53e-07 $l=6.83e-07 $layer=LI1_cond $X=11.562 $Y=1.307
+ $X2=11.562 $Y2=1.99
r99 17 20 7.97992 $w=1.7e-07 $l=2.15346e-07 $layer=LI1_cond $X=11.385 $Y=2.99
+ $X2=11.562 $Y2=2.905
r100 17 18 181.043 $w=1.68e-07 $l=2.775e-06 $layer=LI1_cond $X=11.385 $Y=2.99
+ $X2=8.61 $Y2=2.99
r101 16 18 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=8.39 $Y=2.905
+ $X2=8.61 $Y2=2.99
r102 15 35 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=8.39 $Y=2.1
+ $X2=8.39 $Y2=2.045
r103 15 16 21.0845 $w=4.38e-07 $l=8.05e-07 $layer=LI1_cond $X=8.39 $Y=2.1
+ $X2=8.39 $Y2=2.905
r104 13 29 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.255 $Y=1.21
+ $X2=8.255 $Y2=1.085
r105 13 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.255 $Y=1.21
+ $X2=8.255 $Y2=1.88
r106 4 22 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=11.37
+ $Y=1.84 $X2=11.545 $Y2=1.99
r107 3 35 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=8.3
+ $Y=1.87 $X2=8.445 $Y2=2.045
r108 2 28 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=11.35
+ $Y=0.47 $X2=11.57 $Y2=0.965
r109 2 25 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=11.35
+ $Y=0.47 $X2=11.57 $Y2=0.515
r110 1 32 182 $w=1.7e-07 $l=6.43428e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.47 $X2=8.47 $Y2=1.045
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%A_1849_374# 1 2 3 4 15 18 19 20 21 22 25 27 29
+ 31 36 37 39 47
r109 45 47 10.1363 $w=5.88e-07 $l=5e-07 $layer=LI1_cond $X=9.81 $Y=2.1 $X2=10.31
+ $Y2=2.1
r110 43 45 6.68993 $w=5.88e-07 $l=3.3e-07 $layer=LI1_cond $X=9.48 $Y=2.1
+ $X2=9.81 $Y2=2.1
r111 40 49 7.22832 $w=3.46e-07 $l=2.05e-07 $layer=LI1_cond $X=12.62 $Y=2.035
+ $X2=12.62 $Y2=1.83
r112 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.52 $Y=2.035
+ $X2=12.52 $Y2=2.035
r113 36 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.375 $Y=2.035
+ $X2=12.52 $Y2=2.035
r114 36 37 2.35148 $w=1.4e-07 $l=1.9e-06 $layer=MET1_cond $X=12.375 $Y=2.035
+ $X2=10.475 $Y2=2.035
r115 33 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.33 $Y=2.035
+ $X2=10.33 $Y2=2.035
r116 31 37 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=10.36 $Y=2.035
+ $X2=10.475 $Y2=2.035
r117 31 33 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=10.36 $Y=2.035
+ $X2=10.33 $Y2=2.035
r118 27 40 4.40751 $w=3.46e-07 $l=1.5411e-07 $layer=LI1_cond $X=12.685 $Y=2.16
+ $X2=12.62 $Y2=2.035
r119 27 29 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=12.685 $Y=2.16
+ $X2=12.685 $Y2=2.815
r120 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=12.64 $Y=0.79
+ $X2=12.64 $Y2=0.515
r121 21 49 3.38667 $w=2.2e-07 $l=2.3e-07 $layer=LI1_cond $X=12.39 $Y=1.83
+ $X2=12.62 $Y2=1.83
r122 21 22 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=12.39 $Y=1.83
+ $X2=12.08 $Y2=1.83
r123 19 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.475 $Y=0.875
+ $X2=12.64 $Y2=0.79
r124 19 20 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.475 $Y=0.875
+ $X2=12.08 $Y2=0.875
r125 18 22 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=11.995 $Y=1.72
+ $X2=12.08 $Y2=1.83
r126 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.995 $Y=0.96
+ $X2=12.08 $Y2=0.875
r127 17 18 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=11.995 $Y=0.96
+ $X2=11.995 $Y2=1.72
r128 13 45 4.13774 $w=3.3e-07 $l=2.95e-07 $layer=LI1_cond $X=9.81 $Y=1.805
+ $X2=9.81 $Y2=2.1
r129 13 15 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=9.81 $Y=1.805
+ $X2=9.81 $Y2=1.045
r130 4 40 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.96 $X2=12.685 $Y2=2.135
r131 4 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.96 $X2=12.685 $Y2=2.815
r132 3 47 150 $w=1.7e-07 $l=1.11388e-06 $layer=licon1_PDIFF $count=4 $X=9.245
+ $Y=1.87 $X2=10.31 $Y2=1.97
r133 3 43 300 $w=1.7e-07 $l=2.8058e-07 $layer=licon1_PDIFF $count=2 $X=9.245
+ $Y=1.87 $X2=9.48 $Y2=1.97
r134 2 25 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.495
+ $Y=0.37 $X2=12.64 $Y2=0.515
r135 1 15 182 $w=1.7e-07 $l=6.7611e-07 $layer=licon1_NDIFF $count=1 $X=9.59
+ $Y=0.47 $X2=9.81 $Y2=1.045
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_1%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 42
+ 44 56 70 76 77 80 83 86
r120 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r121 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r122 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 77 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r124 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r125 74 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.14 $Y2=0
r126 74 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.68 $Y2=0
r127 73 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r128 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r129 70 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=13.14 $Y2=0
r130 70 72 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=12.72 $Y2=0
r131 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r132 68 69 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r133 66 69 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=11.76 $Y2=0
r134 66 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r135 65 68 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=11.76
+ $Y2=0
r136 65 66 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r137 63 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=7.91
+ $Y2=0
r138 63 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=8.4
+ $Y2=0
r139 62 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r140 61 62 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r141 58 61 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=7.44
+ $Y2=0
r142 58 59 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r143 56 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.91
+ $Y2=0
r144 56 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r145 55 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r146 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r147 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r148 52 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r149 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r150 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r151 49 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r152 49 51 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r153 47 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r154 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r155 44 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.785
+ $Y2=0
r156 44 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r157 42 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r158 42 59 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=2.64
+ $Y2=0
r159 40 68 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=11.915 $Y=0
+ $X2=11.76 $Y2=0
r160 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.915 $Y=0
+ $X2=12.08 $Y2=0
r161 39 72 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=12.245 $Y=0
+ $X2=12.72 $Y2=0
r162 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.245 $Y=0
+ $X2=12.08 $Y2=0
r163 37 54 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.16
+ $Y2=0
r164 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.34
+ $Y2=0
r165 36 58 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.425 $Y=0
+ $X2=2.64 $Y2=0
r166 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.34
+ $Y2=0
r167 32 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0
r168 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0.515
r169 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.08 $Y=0.085
+ $X2=12.08 $Y2=0
r170 28 30 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.08 $Y=0.085
+ $X2=12.08 $Y2=0.455
r171 24 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r172 24 26 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.365
r173 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.085
+ $X2=2.34 $Y2=0
r174 20 22 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.34 $Y=0.085
+ $X2=2.34 $Y2=0.565
r175 16 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r176 16 18 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.475
r177 5 34 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=12.97
+ $Y=0.37 $X2=13.14 $Y2=0.515
r178 4 30 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=11.86
+ $Y=0.37 $X2=12.08 $Y2=0.455
r179 3 26 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.69
+ $Y=0.37 $X2=7.91 $Y2=0.365
r180 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.2
+ $Y=0.42 $X2=2.34 $Y2=0.565
r181 1 18 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.56 $X2=0.785 $Y2=0.475
.ends

