# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__o221ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o221ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.645000 1.350000 3.975000 1.950000 ;
        RECT 3.645000 1.950000 5.635000 2.120000 ;
        RECT 4.925000 1.350000 5.635000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.350000 4.675000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.350000 2.275000 1.950000 ;
        RECT 1.085000 1.950000 3.405000 2.120000 ;
        RECT 3.075000 1.350000 3.405000 1.950000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.520000 1.350000 2.850000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.232000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.595000 0.875000 2.290000 ;
        RECT 0.605000 2.290000 4.615000 2.460000 ;
        RECT 0.605000 2.460000 0.855000 2.980000 ;
        RECT 2.365000 2.460000 2.695000 2.735000 ;
        RECT 4.365000 2.460000 4.615000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 5.760000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 5.950000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.255000 1.305000 0.425000 ;
      RECT 0.115000  0.425000 0.365000 1.130000 ;
      RECT 0.155000  1.950000 0.405000 3.245000 ;
      RECT 1.055000  0.425000 1.305000 1.010000 ;
      RECT 1.055000  1.010000 3.280000 1.180000 ;
      RECT 1.055000  2.630000 1.695000 3.245000 ;
      RECT 1.535000  0.255000 3.710000 0.425000 ;
      RECT 1.535000  0.425000 1.865000 0.820000 ;
      RECT 1.865000  2.630000 2.195000 2.905000 ;
      RECT 1.865000  2.905000 3.195000 3.075000 ;
      RECT 2.045000  0.595000 2.215000 1.010000 ;
      RECT 2.395000  0.425000 2.725000 0.820000 ;
      RECT 2.865000  2.630000 3.195000 2.905000 ;
      RECT 2.895000  0.595000 3.280000 1.010000 ;
      RECT 3.365000  2.630000 3.695000 3.245000 ;
      RECT 3.460000  0.425000 3.710000 1.010000 ;
      RECT 3.460000  1.010000 5.645000 1.180000 ;
      RECT 3.865000  2.630000 4.195000 2.905000 ;
      RECT 3.865000  2.905000 5.145000 3.075000 ;
      RECT 3.880000  0.085000 4.210000 0.820000 ;
      RECT 4.380000  0.405000 4.710000 1.010000 ;
      RECT 4.815000  2.290000 5.145000 2.905000 ;
      RECT 4.880000  0.085000 5.210000 0.820000 ;
      RECT 5.315000  2.290000 5.645000 3.245000 ;
      RECT 5.390000  0.405000 5.645000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__o221ai_2
END LIBRARY
