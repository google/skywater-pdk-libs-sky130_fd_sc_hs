* File: sky130_fd_sc_hs__einvp_2.pxi.spice
* Created: Tue Sep  1 20:05:03 2020
* 
x_PM_SKY130_FD_SC_HS__EINVP_2%A N_A_c_75_n N_A_M1003_g N_A_c_71_n N_A_M1001_g
+ N_A_c_76_n N_A_M1005_g N_A_c_72_n N_A_M1009_g A N_A_c_74_n
+ PM_SKY130_FD_SC_HS__EINVP_2%A
x_PM_SKY130_FD_SC_HS__EINVP_2%A_263_323# N_A_263_323#_M1000_s
+ N_A_263_323#_M1004_s N_A_263_323#_c_122_n N_A_263_323#_M1006_g
+ N_A_263_323#_c_115_n N_A_263_323#_c_116_n N_A_263_323#_c_125_n
+ N_A_263_323#_M1007_g N_A_263_323#_c_117_n N_A_263_323#_c_118_n
+ N_A_263_323#_c_119_n N_A_263_323#_c_120_n N_A_263_323#_c_121_n
+ PM_SKY130_FD_SC_HS__EINVP_2%A_263_323#
x_PM_SKY130_FD_SC_HS__EINVP_2%TE N_TE_c_176_n N_TE_M1002_g N_TE_c_177_n
+ N_TE_c_178_n N_TE_c_179_n N_TE_M1008_g N_TE_c_180_n N_TE_c_181_n N_TE_M1000_g
+ N_TE_c_188_n N_TE_M1004_g N_TE_c_183_n N_TE_c_184_n N_TE_c_190_n N_TE_c_185_n
+ TE N_TE_c_186_n N_TE_c_187_n PM_SKY130_FD_SC_HS__EINVP_2%TE
x_PM_SKY130_FD_SC_HS__EINVP_2%A_27_368# N_A_27_368#_M1003_d N_A_27_368#_M1005_d
+ N_A_27_368#_M1007_s N_A_27_368#_c_243_n N_A_27_368#_c_244_n
+ N_A_27_368#_c_245_n N_A_27_368#_c_246_n N_A_27_368#_c_241_n
+ N_A_27_368#_c_242_n N_A_27_368#_c_247_n PM_SKY130_FD_SC_HS__EINVP_2%A_27_368#
x_PM_SKY130_FD_SC_HS__EINVP_2%Z N_Z_M1001_s N_Z_M1003_s N_Z_c_291_n Z Z Z Z Z
+ PM_SKY130_FD_SC_HS__EINVP_2%Z
x_PM_SKY130_FD_SC_HS__EINVP_2%VPWR N_VPWR_M1006_d N_VPWR_M1004_d N_VPWR_c_314_n
+ N_VPWR_c_315_n N_VPWR_c_316_n VPWR N_VPWR_c_317_n N_VPWR_c_318_n
+ N_VPWR_c_319_n N_VPWR_c_313_n PM_SKY130_FD_SC_HS__EINVP_2%VPWR
x_PM_SKY130_FD_SC_HS__EINVP_2%A_36_74# N_A_36_74#_M1001_d N_A_36_74#_M1009_d
+ N_A_36_74#_M1008_s N_A_36_74#_c_349_n N_A_36_74#_c_350_n N_A_36_74#_c_351_n
+ N_A_36_74#_c_352_n N_A_36_74#_c_353_n N_A_36_74#_c_354_n N_A_36_74#_c_355_n
+ PM_SKY130_FD_SC_HS__EINVP_2%A_36_74#
x_PM_SKY130_FD_SC_HS__EINVP_2%VGND N_VGND_M1002_d N_VGND_M1000_d N_VGND_c_397_n
+ N_VGND_c_398_n N_VGND_c_399_n VGND N_VGND_c_400_n N_VGND_c_401_n
+ N_VGND_c_402_n N_VGND_c_403_n PM_SKY130_FD_SC_HS__EINVP_2%VGND
cc_1 VNB N_A_c_71_n 0.0203982f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.22
cc_2 VNB N_A_c_72_n 0.0159117f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.22
cc_3 VNB A 0.0113831f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_74_n 0.10253f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.492
cc_5 VNB N_A_263_323#_c_115_n 0.00539409f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.22
cc_6 VNB N_A_263_323#_c_116_n 0.00376765f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_7 VNB N_A_263_323#_c_117_n 0.00269832f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_8 VNB N_A_263_323#_c_118_n 0.0160163f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.492
cc_9 VNB N_A_263_323#_c_119_n 0.0164879f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.492
cc_10 VNB N_A_263_323#_c_120_n 0.00526886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_263_323#_c_121_n 0.0101994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_TE_c_176_n 0.0145546f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_13 VNB N_TE_c_177_n 0.0126145f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.22
cc_14 VNB N_TE_c_178_n 0.00751923f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_15 VNB N_TE_c_179_n 0.0161538f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_16 VNB N_TE_c_180_n 0.026203f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_17 VNB N_TE_c_181_n 0.0333291f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_18 VNB N_TE_M1000_g 0.0120118f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_19 VNB N_TE_c_183_n 0.0251423f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.492
cc_20 VNB N_TE_c_184_n 0.00535066f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_21 VNB N_TE_c_185_n 0.0342067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_TE_c_186_n 0.0588596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_TE_c_187_n 0.00566583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_368#_c_241_n 0.00845447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_368#_c_242_n 0.00299021f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_26 VNB N_Z_c_291_n 6.47547e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_27 VNB Z 0.0033102f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_28 VNB N_VPWR_c_313_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_36_74#_c_349_n 0.0222939f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_30 VNB N_A_36_74#_c_350_n 0.00449328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_36_74#_c_351_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.492
cc_32 VNB N_A_36_74#_c_352_n 4.66303e-19 $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.492
cc_33 VNB N_A_36_74#_c_353_n 0.00668482f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.492
cc_34 VNB N_A_36_74#_c_354_n 0.00289968f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.492
cc_35 VNB N_A_36_74#_c_355_n 0.00892448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_397_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_37 VNB N_VGND_c_398_n 0.0109649f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_38 VNB N_VGND_c_399_n 0.0418368f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_39 VNB N_VGND_c_400_n 0.0374035f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_40 VNB N_VGND_c_401_n 0.0327804f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_41 VNB N_VGND_c_402_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_403_n 0.215736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A_c_75_n 0.0184183f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_44 VPB N_A_c_76_n 0.0145627f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_45 VPB N_A_c_74_n 0.0169982f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.492
cc_46 VPB N_A_263_323#_c_122_n 0.0152711f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_47 VPB N_A_263_323#_c_115_n 0.00587316f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.22
cc_48 VPB N_A_263_323#_c_116_n 0.00457213f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=0.74
cc_49 VPB N_A_263_323#_c_125_n 0.0191108f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=0.74
cc_50 VPB N_A_263_323#_c_117_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_51 VPB N_A_263_323#_c_118_n 0.0237004f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.492
cc_52 VPB N_A_263_323#_c_119_n 0.0242617f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.492
cc_53 VPB N_A_263_323#_c_121_n 0.0238269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_TE_c_188_n 0.0221231f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_55 VPB N_TE_c_183_n 0.0347972f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.492
cc_56 VPB N_TE_c_190_n 0.0343249f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_57 VPB N_A_27_368#_c_243_n 0.0419775f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=0.74
cc_58 VPB N_A_27_368#_c_244_n 0.00522128f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_59 VPB N_A_27_368#_c_245_n 0.00935849f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_60 VPB N_A_27_368#_c_246_n 0.00282099f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.492
cc_61 VPB N_A_27_368#_c_247_n 0.00275579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB Z 0.00200122f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=0.74
cc_63 VPB N_VPWR_c_314_n 0.00739602f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_64 VPB N_VPWR_c_315_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_65 VPB N_VPWR_c_316_n 0.0418872f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.492
cc_66 VPB N_VPWR_c_317_n 0.0375082f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.492
cc_67 VPB N_VPWR_c_318_n 0.0334651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_319_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_313_n 0.0730506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 N_A_c_76_n N_A_263_323#_c_122_n 0.0087792f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A_c_74_n N_A_263_323#_c_116_n 0.00635824f $X=0.955 $Y=1.492 $X2=0 $Y2=0
cc_72 N_A_c_72_n N_TE_c_176_n 0.00855951f $X=0.97 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_73 N_A_c_74_n N_TE_c_178_n 0.00855951f $X=0.955 $Y=1.492 $X2=0 $Y2=0
cc_74 N_A_c_75_n N_A_27_368#_c_243_n 0.00863263f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_75 A N_A_27_368#_c_243_n 0.0149782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_c_74_n N_A_27_368#_c_243_n 0.00185549f $X=0.955 $Y=1.492 $X2=0 $Y2=0
cc_77 N_A_c_75_n N_A_27_368#_c_244_n 0.0140817f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_78 N_A_c_76_n N_A_27_368#_c_244_n 0.0117394f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_c_76_n N_A_27_368#_c_246_n 0.00653858f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_74_n N_A_27_368#_c_246_n 8.22435e-19 $X=0.955 $Y=1.492 $X2=0 $Y2=0
cc_81 N_A_c_74_n N_A_27_368#_c_242_n 0.00406866f $X=0.955 $Y=1.492 $X2=0 $Y2=0
cc_82 N_A_c_71_n N_Z_c_291_n 0.00215527f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_83 N_A_c_72_n N_Z_c_291_n 0.00757448f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_84 N_A_c_75_n Z 0.00265652f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_c_71_n Z 0.00131177f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_86 N_A_c_76_n Z 0.0142908f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_c_72_n Z 8.7164e-19 $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_88 A Z 0.0277568f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A_c_74_n Z 0.0377983f $X=0.955 $Y=1.492 $X2=0 $Y2=0
cc_90 N_A_c_75_n N_VPWR_c_317_n 0.00278271f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_c_76_n N_VPWR_c_317_n 0.00278271f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_c_75_n N_VPWR_c_313_n 0.00357317f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_c_76_n N_VPWR_c_313_n 0.00353907f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_c_71_n N_A_36_74#_c_349_n 0.00929919f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_95 N_A_c_72_n N_A_36_74#_c_349_n 6.05004e-19 $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_96 A N_A_36_74#_c_349_n 0.0228393f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A_c_74_n N_A_36_74#_c_349_n 0.00186453f $X=0.955 $Y=1.492 $X2=0 $Y2=0
cc_98 N_A_c_71_n N_A_36_74#_c_350_n 0.0100245f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_99 N_A_c_72_n N_A_36_74#_c_350_n 0.0120332f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_100 N_A_c_71_n N_A_36_74#_c_351_n 0.00282152f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A_c_72_n N_A_36_74#_c_352_n 4.60747e-19 $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_102 N_A_c_72_n N_A_36_74#_c_354_n 0.0015676f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_103 N_A_c_71_n N_VGND_c_400_n 0.00278247f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_104 N_A_c_72_n N_VGND_c_400_n 0.00278271f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_105 N_A_c_71_n N_VGND_c_403_n 0.00357229f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A_c_72_n N_VGND_c_403_n 0.00353526f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A_263_323#_c_115_n N_TE_c_177_n 0.012678f $X=1.78 $Y=1.69 $X2=0 $Y2=0
cc_108 N_A_263_323#_c_116_n N_TE_c_178_n 0.012678f $X=1.48 $Y=1.69 $X2=0 $Y2=0
cc_109 N_A_263_323#_c_118_n N_TE_c_180_n 0.00297448f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_110 N_A_263_323#_c_121_n N_TE_c_180_n 0.012678f $X=2.415 $Y=1.72 $X2=0 $Y2=0
cc_111 N_A_263_323#_c_120_n N_TE_c_181_n 0.00297448f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_112 N_A_263_323#_c_118_n N_TE_M1000_g 0.00628076f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_113 N_A_263_323#_c_120_n N_TE_M1000_g 0.00915681f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_114 N_A_263_323#_c_118_n N_TE_c_188_n 0.00325651f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_115 N_A_263_323#_c_118_n N_TE_c_183_n 0.0103964f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_116 N_A_263_323#_c_119_n N_TE_c_183_n 0.0190575f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_117 N_A_263_323#_c_117_n N_TE_c_184_n 0.012678f $X=1.855 $Y=1.69 $X2=0 $Y2=0
cc_118 N_A_263_323#_c_118_n N_TE_c_190_n 0.00723932f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_119 N_A_263_323#_c_120_n N_TE_c_186_n 0.00115908f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_120 N_A_263_323#_c_120_n N_TE_c_187_n 0.0247075f $X=2.635 $Y=0.95 $X2=0 $Y2=0
cc_121 N_A_263_323#_c_122_n N_A_27_368#_c_244_n 0.00125031f $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_122 N_A_263_323#_c_122_n N_A_27_368#_c_246_n 0.00442794f $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_123 N_A_263_323#_c_116_n N_A_27_368#_c_246_n 0.00167013f $X=1.48 $Y=1.69
+ $X2=0 $Y2=0
cc_124 N_A_263_323#_c_115_n N_A_27_368#_c_241_n 0.00844732f $X=1.78 $Y=1.69
+ $X2=0 $Y2=0
cc_125 N_A_263_323#_c_116_n N_A_27_368#_c_241_n 0.00885948f $X=1.48 $Y=1.69
+ $X2=0 $Y2=0
cc_126 N_A_263_323#_c_117_n N_A_27_368#_c_241_n 0.00745155f $X=1.855 $Y=1.69
+ $X2=0 $Y2=0
cc_127 N_A_263_323#_c_118_n N_A_27_368#_c_241_n 0.0109091f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_128 N_A_263_323#_c_119_n N_A_27_368#_c_241_n 0.00133801f $X=2.58 $Y=1.72
+ $X2=0 $Y2=0
cc_129 N_A_263_323#_c_121_n N_A_27_368#_c_241_n 0.00304417f $X=2.415 $Y=1.72
+ $X2=0 $Y2=0
cc_130 N_A_263_323#_c_122_n N_A_27_368#_c_247_n 5.59846e-19 $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_131 N_A_263_323#_c_125_n N_A_27_368#_c_247_n 0.015206f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_132 N_A_263_323#_c_117_n N_A_27_368#_c_247_n 0.00315233f $X=1.855 $Y=1.69
+ $X2=0 $Y2=0
cc_133 N_A_263_323#_c_118_n N_A_27_368#_c_247_n 0.0796672f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_134 N_A_263_323#_c_119_n N_A_27_368#_c_247_n 0.00101418f $X=2.58 $Y=1.72
+ $X2=0 $Y2=0
cc_135 N_A_263_323#_c_121_n N_A_27_368#_c_247_n 0.0100643f $X=2.415 $Y=1.72
+ $X2=0 $Y2=0
cc_136 N_A_263_323#_c_122_n N_VPWR_c_314_n 0.0154116f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_263_323#_c_115_n N_VPWR_c_314_n 0.00276433f $X=1.78 $Y=1.69 $X2=0
+ $Y2=0
cc_138 N_A_263_323#_c_125_n N_VPWR_c_314_n 0.00718907f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_263_323#_c_118_n N_VPWR_c_316_n 0.0270962f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_140 N_A_263_323#_c_122_n N_VPWR_c_317_n 0.00413917f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A_263_323#_c_125_n N_VPWR_c_318_n 0.00445602f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_263_323#_c_118_n N_VPWR_c_318_n 0.0146357f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_143 N_A_263_323#_c_122_n N_VPWR_c_313_n 0.0081781f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_A_263_323#_c_125_n N_VPWR_c_313_n 0.00862391f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_A_263_323#_c_118_n N_VPWR_c_313_n 0.0121141f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_146 N_A_263_323#_c_116_n N_A_36_74#_c_353_n 6.578e-19 $X=1.48 $Y=1.69 $X2=0
+ $Y2=0
cc_147 N_A_263_323#_c_118_n N_A_36_74#_c_353_n 0.0125516f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_148 N_A_263_323#_c_121_n N_A_36_74#_c_353_n 4.74394e-19 $X=2.415 $Y=1.72
+ $X2=0 $Y2=0
cc_149 N_A_263_323#_c_120_n N_A_36_74#_c_355_n 0.0217181f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_150 N_A_263_323#_c_120_n N_VGND_c_403_n 0.0031213f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_151 N_TE_c_178_n N_A_27_368#_c_241_n 0.00415283f $X=1.475 $Y=1.26 $X2=0 $Y2=0
cc_152 N_TE_c_180_n N_A_27_368#_c_241_n 0.00179693f $X=2.265 $Y=1.26 $X2=0 $Y2=0
cc_153 N_TE_c_176_n N_Z_c_291_n 2.18758e-19 $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_154 N_TE_c_178_n Z 2.10146e-19 $X=1.475 $Y=1.26 $X2=0 $Y2=0
cc_155 N_TE_c_188_n N_VPWR_c_316_n 0.0152974f $X=2.855 $Y=2.245 $X2=0 $Y2=0
cc_156 N_TE_c_190_n N_VPWR_c_316_n 0.010791f $X=3.06 $Y=2.17 $X2=0 $Y2=0
cc_157 N_TE_c_188_n N_VPWR_c_318_n 0.00413917f $X=2.855 $Y=2.245 $X2=0 $Y2=0
cc_158 N_TE_c_188_n N_VPWR_c_313_n 0.00822528f $X=2.855 $Y=2.245 $X2=0 $Y2=0
cc_159 N_TE_c_176_n N_A_36_74#_c_350_n 9.48753e-19 $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_160 N_TE_c_176_n N_A_36_74#_c_352_n 9.29165e-19 $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_161 N_TE_c_176_n N_A_36_74#_c_353_n 0.00741157f $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_162 N_TE_c_177_n N_A_36_74#_c_353_n 0.00615573f $X=1.755 $Y=1.26 $X2=0 $Y2=0
cc_163 N_TE_c_178_n N_A_36_74#_c_353_n 0.00364399f $X=1.475 $Y=1.26 $X2=0 $Y2=0
cc_164 N_TE_c_179_n N_A_36_74#_c_353_n 0.00753496f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_165 N_TE_c_180_n N_A_36_74#_c_353_n 0.0112425f $X=2.265 $Y=1.26 $X2=0 $Y2=0
cc_166 N_TE_c_181_n N_A_36_74#_c_353_n 4.36766e-19 $X=2.34 $Y=1.185 $X2=0 $Y2=0
cc_167 N_TE_c_184_n N_A_36_74#_c_353_n 0.00251882f $X=1.83 $Y=1.26 $X2=0 $Y2=0
cc_168 N_TE_c_179_n N_A_36_74#_c_355_n 0.00130964f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_169 N_TE_c_186_n N_A_36_74#_c_355_n 0.0106764f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_170 N_TE_c_187_n N_A_36_74#_c_355_n 0.0179335f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_171 N_TE_c_176_n N_VGND_c_397_n 0.0100283f $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_172 N_TE_c_177_n N_VGND_c_397_n 7.11061e-19 $X=1.755 $Y=1.26 $X2=0 $Y2=0
cc_173 N_TE_c_179_n N_VGND_c_397_n 0.0134095f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_174 N_TE_c_185_n N_VGND_c_399_n 0.00727925f $X=3.06 $Y=1.27 $X2=0 $Y2=0
cc_175 N_TE_c_186_n N_VGND_c_399_n 0.0124285f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_176 N_TE_c_187_n N_VGND_c_399_n 0.0318479f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_177 N_TE_c_176_n N_VGND_c_400_n 0.00383152f $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_178 N_TE_c_179_n N_VGND_c_401_n 0.00383152f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_179 N_TE_c_186_n N_VGND_c_401_n 0.0128697f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_180 N_TE_c_187_n N_VGND_c_401_n 0.0208821f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_181 N_TE_c_176_n N_VGND_c_403_n 0.00757637f $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_182 N_TE_c_179_n N_VGND_c_403_n 0.00762539f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_183 N_TE_c_186_n N_VGND_c_403_n 0.011158f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_184 N_TE_c_187_n N_VGND_c_403_n 0.0123609f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_185 N_A_27_368#_c_244_n N_Z_M1003_s 0.00197722f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_186 N_A_27_368#_c_243_n Z 0.0279378f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_27_368#_c_244_n Z 0.0168986f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_188 N_A_27_368#_c_246_n Z 0.0782308f $X=1.18 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_27_368#_c_242_n Z 0.01398f $X=1.265 $Y=1.565 $X2=0 $Y2=0
cc_190 N_A_27_368#_c_244_n N_VPWR_c_314_n 0.0123543f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_191 N_A_27_368#_c_246_n N_VPWR_c_314_n 0.0691797f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_27_368#_c_241_n N_VPWR_c_314_n 0.0199131f $X=1.915 $Y=1.565 $X2=0
+ $Y2=0
cc_193 N_A_27_368#_c_247_n N_VPWR_c_314_n 0.0762465f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_27_368#_c_244_n N_VPWR_c_317_n 0.0582081f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_195 N_A_27_368#_c_245_n N_VPWR_c_317_n 0.0179217f $X=0.365 $Y=2.99 $X2=0
+ $Y2=0
cc_196 N_A_27_368#_c_247_n N_VPWR_c_318_n 0.0110241f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_197 N_A_27_368#_c_244_n N_VPWR_c_313_n 0.0326718f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_198 N_A_27_368#_c_245_n N_VPWR_c_313_n 0.00971942f $X=0.365 $Y=2.99 $X2=0
+ $Y2=0
cc_199 N_A_27_368#_c_247_n N_VPWR_c_313_n 0.00909194f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_27_368#_c_241_n N_A_36_74#_c_353_n 0.0681198f $X=1.915 $Y=1.565 $X2=0
+ $Y2=0
cc_201 N_A_27_368#_c_241_n N_A_36_74#_c_354_n 3.84494e-19 $X=1.915 $Y=1.565
+ $X2=0 $Y2=0
cc_202 N_A_27_368#_c_242_n N_A_36_74#_c_354_n 0.0154601f $X=1.265 $Y=1.565 $X2=0
+ $Y2=0
cc_203 N_Z_M1001_s N_A_36_74#_c_350_n 0.00189202f $X=0.615 $Y=0.37 $X2=0 $Y2=0
cc_204 N_Z_c_291_n N_A_36_74#_c_350_n 0.0124268f $X=0.755 $Y=0.82 $X2=0 $Y2=0
cc_205 N_Z_c_291_n N_A_36_74#_c_352_n 0.0187012f $X=0.755 $Y=0.82 $X2=0 $Y2=0
cc_206 N_Z_c_291_n N_A_36_74#_c_354_n 0.0135667f $X=0.755 $Y=0.82 $X2=0 $Y2=0
cc_207 N_A_36_74#_c_350_n N_VGND_c_397_n 0.0112234f $X=1.1 $Y=0.34 $X2=0 $Y2=0
cc_208 N_A_36_74#_c_353_n N_VGND_c_397_n 0.0216086f $X=1.95 $Y=1.225 $X2=0 $Y2=0
cc_209 N_A_36_74#_c_355_n N_VGND_c_397_n 0.0240263f $X=2.045 $Y=0.515 $X2=0
+ $Y2=0
cc_210 N_A_36_74#_c_350_n N_VGND_c_400_n 0.050626f $X=1.1 $Y=0.34 $X2=0 $Y2=0
cc_211 N_A_36_74#_c_351_n N_VGND_c_400_n 0.0235688f $X=0.49 $Y=0.34 $X2=0 $Y2=0
cc_212 N_A_36_74#_c_355_n N_VGND_c_401_n 0.0115122f $X=2.045 $Y=0.515 $X2=0
+ $Y2=0
cc_213 N_A_36_74#_c_350_n N_VGND_c_403_n 0.028285f $X=1.1 $Y=0.34 $X2=0 $Y2=0
cc_214 N_A_36_74#_c_351_n N_VGND_c_403_n 0.0127152f $X=0.49 $Y=0.34 $X2=0 $Y2=0
cc_215 N_A_36_74#_c_355_n N_VGND_c_403_n 0.0095288f $X=2.045 $Y=0.515 $X2=0
+ $Y2=0
