* File: sky130_fd_sc_hs__o221a_2.pxi.spice
* Created: Thu Aug 27 20:59:18 2020
* 
x_PM_SKY130_FD_SC_HS__O221A_2%C1 N_C1_c_84_n N_C1_M1013_g N_C1_c_81_n
+ N_C1_M1006_g C1 N_C1_c_83_n PM_SKY130_FD_SC_HS__O221A_2%C1
x_PM_SKY130_FD_SC_HS__O221A_2%B1 N_B1_M1010_g N_B1_c_112_n N_B1_M1002_g B1
+ N_B1_c_110_n N_B1_c_111_n PM_SKY130_FD_SC_HS__O221A_2%B1
x_PM_SKY130_FD_SC_HS__O221A_2%B2 N_B2_c_148_n N_B2_M1003_g N_B2_c_149_n
+ N_B2_c_150_n N_B2_c_151_n N_B2_M1008_g B2 B2 PM_SKY130_FD_SC_HS__O221A_2%B2
x_PM_SKY130_FD_SC_HS__O221A_2%A2 N_A2_c_187_n N_A2_M1011_g N_A2_M1012_g A2
+ N_A2_c_189_n PM_SKY130_FD_SC_HS__O221A_2%A2
x_PM_SKY130_FD_SC_HS__O221A_2%A1 N_A1_c_216_n N_A1_M1009_g N_A1_M1004_g A1
+ N_A1_c_218_n PM_SKY130_FD_SC_HS__O221A_2%A1
x_PM_SKY130_FD_SC_HS__O221A_2%A_27_368# N_A_27_368#_M1006_s N_A_27_368#_M1013_s
+ N_A_27_368#_M1008_d N_A_27_368#_M1000_g N_A_27_368#_c_252_n
+ N_A_27_368#_M1001_g N_A_27_368#_c_253_n N_A_27_368#_M1007_g
+ N_A_27_368#_c_255_n N_A_27_368#_c_264_n N_A_27_368#_M1005_g
+ N_A_27_368#_c_256_n N_A_27_368#_c_265_n N_A_27_368#_c_257_n
+ N_A_27_368#_c_258_n N_A_27_368#_c_276_n N_A_27_368#_c_267_n
+ N_A_27_368#_c_296_n N_A_27_368#_c_259_n N_A_27_368#_c_269_n
+ N_A_27_368#_c_260_n N_A_27_368#_c_293_n N_A_27_368#_c_261_n
+ PM_SKY130_FD_SC_HS__O221A_2%A_27_368#
x_PM_SKY130_FD_SC_HS__O221A_2%VPWR N_VPWR_M1013_d N_VPWR_M1009_d N_VPWR_M1005_s
+ N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n VPWR
+ N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_372_n
+ N_VPWR_c_363_n PM_SKY130_FD_SC_HS__O221A_2%VPWR
x_PM_SKY130_FD_SC_HS__O221A_2%X N_X_M1000_s N_X_M1001_d N_X_c_415_n N_X_c_416_n
+ N_X_c_412_n X X N_X_c_413_n X PM_SKY130_FD_SC_HS__O221A_2%X
x_PM_SKY130_FD_SC_HS__O221A_2%A_165_74# N_A_165_74#_M1006_d N_A_165_74#_M1003_d
+ N_A_165_74#_c_448_n N_A_165_74#_c_449_n N_A_165_74#_c_450_n
+ PM_SKY130_FD_SC_HS__O221A_2%A_165_74#
x_PM_SKY130_FD_SC_HS__O221A_2%A_264_74# N_A_264_74#_M1010_d N_A_264_74#_M1012_d
+ N_A_264_74#_c_474_n N_A_264_74#_c_475_n N_A_264_74#_c_476_n
+ PM_SKY130_FD_SC_HS__O221A_2%A_264_74#
x_PM_SKY130_FD_SC_HS__O221A_2%VGND N_VGND_M1012_s N_VGND_M1004_d N_VGND_M1007_d
+ N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n N_VGND_c_513_n
+ N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n VGND N_VGND_c_517_n
+ N_VGND_c_518_n PM_SKY130_FD_SC_HS__O221A_2%VGND
cc_1 VNB N_C1_c_81_n 0.0227378f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.22
cc_2 VNB C1 0.0159976f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_C1_c_83_n 0.0913524f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_4 VNB N_B1_M1010_g 0.0263143f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_5 VNB N_B1_c_110_n 0.00333483f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_6 VNB N_B1_c_111_n 0.0396956f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.492
cc_7 VNB N_B2_c_148_n 0.0181556f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_8 VNB N_B2_c_149_n 0.0318136f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.22
cc_9 VNB N_B2_c_150_n 0.0122502f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.74
cc_10 VNB N_B2_c_151_n 0.00898421f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.74
cc_11 VNB B2 0.00636131f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_12 VNB N_A2_c_187_n 0.0269958f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_13 VNB N_A2_M1012_g 0.027284f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.74
cc_14 VNB N_A2_c_189_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_15 VNB N_A1_c_216_n 0.0247514f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_16 VNB N_A1_M1004_g 0.0261039f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.74
cc_17 VNB N_A1_c_218_n 0.00552033f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_18 VNB N_A_27_368#_M1000_g 0.0241917f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_19 VNB N_A_27_368#_c_252_n 0.0278552f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_20 VNB N_A_27_368#_c_253_n 0.00638712f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_21 VNB N_A_27_368#_M1007_g 0.0251809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_368#_c_255_n 0.0150953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_368#_c_256_n 0.0206399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_368#_c_257_n 0.0204696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_368#_c_258_n 0.00460576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_368#_c_259_n 2.18704e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_368#_c_260_n 0.00797994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_368#_c_261_n 0.00257315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_363_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_412_n 0.00795141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_413_n 0.00274256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB X 0.00577223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_165_74#_c_448_n 0.00342538f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.492
cc_34 VNB N_A_165_74#_c_449_n 0.00716791f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_35 VNB N_A_165_74#_c_450_n 0.00704577f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.492
cc_36 VNB N_A_264_74#_c_474_n 0.0300192f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_37 VNB N_A_264_74#_c_475_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_38 VNB N_A_264_74#_c_476_n 0.00313103f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_39 VNB N_VGND_c_509_n 0.0106116f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_40 VNB N_VGND_c_510_n 0.017767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_511_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_512_n 0.0506881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_513_n 0.0648512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_514_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_515_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_516_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_517_n 0.0221763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_518_n 0.299576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VPB N_C1_c_84_n 0.0206815f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_50 VPB N_C1_c_83_n 0.010241f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_51 VPB N_B1_c_112_n 0.0180105f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=0.74
cc_52 VPB N_B1_c_110_n 0.00384845f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_53 VPB N_B1_c_111_n 0.0212207f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.492
cc_54 VPB N_B2_c_151_n 0.0262824f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=0.74
cc_55 VPB B2 0.00513457f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_56 VPB N_A2_c_187_n 0.0285966f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_57 VPB N_A2_c_189_n 0.00241345f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_58 VPB N_A1_c_216_n 0.0290501f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_59 VPB N_A1_c_218_n 0.00363387f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_60 VPB N_A_27_368#_c_252_n 0.0242205f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_61 VPB N_A_27_368#_c_255_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_368#_c_264_n 0.0257687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_368#_c_265_n 0.0315121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_368#_c_258_n 0.00446037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_27_368#_c_267_n 0.00358314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_27_368#_c_259_n 0.00290198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_368#_c_269_n 0.0161978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_364_n 0.02606f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_69 VPB N_VPWR_c_365_n 0.0143582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_366_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_367_n 0.0644986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_368_n 0.0196898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_369_n 0.0577377f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_370_n 0.0194151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_371_n 0.0174777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_372_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_363_n 0.112271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_X_c_415_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.492
cc_79 VPB N_X_c_416_n 0.00472837f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_80 VPB N_X_c_412_n 8.52106e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 N_C1_c_81_n N_B1_M1010_g 0.024596f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_82 N_C1_c_83_n N_B1_c_110_n 8.785e-19 $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_83 N_C1_c_83_n N_B1_c_111_n 0.0144443f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_84 N_C1_c_84_n N_A_27_368#_c_265_n 0.0135071f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_85 N_C1_c_81_n N_A_27_368#_c_257_n 0.00869286f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_86 N_C1_c_84_n N_A_27_368#_c_258_n 0.00218667f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_87 N_C1_c_81_n N_A_27_368#_c_258_n 0.00554011f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_88 C1 N_A_27_368#_c_258_n 0.0267371f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_C1_c_83_n N_A_27_368#_c_258_n 0.0248849f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_90 N_C1_c_83_n N_A_27_368#_c_276_n 0.00161321f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_91 N_C1_c_84_n N_A_27_368#_c_269_n 0.0240449f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_92 C1 N_A_27_368#_c_269_n 0.0179404f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_93 N_C1_c_83_n N_A_27_368#_c_269_n 0.00421605f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_94 N_C1_c_81_n N_A_27_368#_c_260_n 0.00306847f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_95 C1 N_A_27_368#_c_260_n 0.00555399f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_96 N_C1_c_83_n N_A_27_368#_c_260_n 0.00823071f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_97 N_C1_c_84_n N_VPWR_c_364_n 0.0164733f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_98 N_C1_c_84_n N_VPWR_c_368_n 0.00481995f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_99 N_C1_c_84_n N_VPWR_c_363_n 0.00508379f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_100 N_C1_c_81_n N_A_165_74#_c_449_n 0.005506f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_101 N_C1_c_81_n N_A_264_74#_c_476_n 2.32508e-19 $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_102 N_C1_c_81_n N_VGND_c_513_n 0.00349296f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_103 N_C1_c_81_n N_VGND_c_518_n 0.00551056f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_104 N_B1_M1010_g N_B2_c_148_n 0.027221f $X=1.245 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_105 N_B1_M1010_g N_B2_c_150_n 3.78334e-19 $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_106 N_B1_c_110_n N_B2_c_150_n 2.50985e-19 $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_107 N_B1_c_111_n N_B2_c_150_n 0.00382197f $X=1.245 $Y=1.557 $X2=0 $Y2=0
cc_108 N_B1_c_112_n N_B2_c_151_n 0.0550619f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_109 N_B1_c_111_n N_B2_c_151_n 0.0104555f $X=1.245 $Y=1.557 $X2=0 $Y2=0
cc_110 N_B1_c_112_n B2 0.00170156f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B1_c_110_n B2 0.0354777f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_112 N_B1_c_111_n B2 0.0108616f $X=1.245 $Y=1.557 $X2=0 $Y2=0
cc_113 N_B1_M1010_g N_A_27_368#_c_257_n 0.00133362f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B1_c_110_n N_A_27_368#_c_258_n 0.0211588f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_115 N_B1_c_111_n N_A_27_368#_c_258_n 0.00217035f $X=1.245 $Y=1.557 $X2=0
+ $Y2=0
cc_116 N_B1_c_112_n N_A_27_368#_c_276_n 0.018068f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_117 N_B1_c_110_n N_A_27_368#_c_276_n 0.0262472f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B1_c_111_n N_A_27_368#_c_276_n 0.00455162f $X=1.245 $Y=1.557 $X2=0
+ $Y2=0
cc_119 N_B1_c_112_n N_A_27_368#_c_267_n 0.00245895f $X=1.585 $Y=1.765 $X2=0
+ $Y2=0
cc_120 N_B1_c_112_n N_VPWR_c_364_n 0.0153074f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_121 N_B1_c_112_n N_VPWR_c_369_n 0.00443511f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B1_c_112_n N_VPWR_c_363_n 0.00460931f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B1_M1010_g N_A_165_74#_c_448_n 0.0123547f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_124 N_B1_M1010_g N_A_165_74#_c_449_n 4.59233e-19 $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_125 N_B1_c_110_n N_A_165_74#_c_449_n 0.00341112f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_126 N_B1_c_111_n N_A_165_74#_c_449_n 3.67352e-19 $X=1.245 $Y=1.557 $X2=0
+ $Y2=0
cc_127 N_B1_M1010_g N_A_165_74#_c_450_n 0.00133243f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_128 N_B1_c_111_n N_A_264_74#_c_474_n 2.29618e-19 $X=1.245 $Y=1.557 $X2=0
+ $Y2=0
cc_129 N_B1_M1010_g N_A_264_74#_c_476_n 0.00591218f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_130 N_B1_c_110_n N_A_264_74#_c_476_n 0.00797323f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_131 N_B1_c_111_n N_A_264_74#_c_476_n 0.00618712f $X=1.245 $Y=1.557 $X2=0
+ $Y2=0
cc_132 N_B1_M1010_g N_VGND_c_513_n 0.00291649f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_133 N_B1_M1010_g N_VGND_c_518_n 0.00360544f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_134 N_B2_c_150_n N_A2_c_187_n 0.0174954f $X=2.08 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_135 N_B2_c_151_n N_A2_c_187_n 0.0200679f $X=2.005 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_136 B2 N_A2_c_187_n 0.00290196f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_137 N_B2_c_149_n N_A2_M1012_g 0.00639049f $X=2.08 $Y=1.335 $X2=0 $Y2=0
cc_138 N_B2_c_150_n N_A2_c_189_n 3.95877e-19 $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_139 B2 N_A2_c_189_n 0.0309799f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_140 N_B2_c_151_n N_A_27_368#_c_276_n 0.0117808f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_141 B2 N_A_27_368#_c_276_n 0.0341134f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_142 N_B2_c_151_n N_A_27_368#_c_267_n 0.0129952f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_143 N_B2_c_151_n N_A_27_368#_c_293_n 0.0012408f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_144 B2 N_A_27_368#_c_293_n 0.0158578f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_145 N_B2_c_151_n N_VPWR_c_364_n 0.00215867f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_146 N_B2_c_151_n N_VPWR_c_369_n 0.00481995f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_147 N_B2_c_151_n N_VPWR_c_363_n 0.00508379f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_148 N_B2_c_148_n N_A_165_74#_c_448_n 0.00917015f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_149 N_B2_c_148_n N_A_165_74#_c_450_n 0.0096459f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_150 N_B2_c_148_n N_A_264_74#_c_474_n 0.0116015f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_151 N_B2_c_149_n N_A_264_74#_c_474_n 0.0122779f $X=2.08 $Y=1.335 $X2=0 $Y2=0
cc_152 B2 N_A_264_74#_c_474_n 0.0510553f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_153 B2 N_A_264_74#_c_476_n 0.00465791f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_154 N_B2_c_148_n N_VGND_c_509_n 0.00383008f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_155 N_B2_c_148_n N_VGND_c_513_n 0.00292759f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_156 N_B2_c_148_n N_VGND_c_518_n 0.00363909f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_157 N_A2_c_187_n N_A1_c_216_n 0.0574184f $X=2.575 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A2_c_189_n N_A1_c_216_n 7.2702e-19 $X=2.65 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A2_M1012_g N_A1_M1004_g 0.0195038f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_c_187_n N_A1_c_218_n 0.00231456f $X=2.575 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A2_c_189_n N_A1_c_218_n 0.0320816f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A2_c_187_n N_A_27_368#_c_267_n 0.0200073f $X=2.575 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A2_c_187_n N_A_27_368#_c_296_n 0.0170894f $X=2.575 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A2_c_189_n N_A_27_368#_c_296_n 0.0226548f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A2_c_187_n N_VPWR_c_369_n 0.0049405f $X=2.575 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A2_c_187_n N_VPWR_c_363_n 0.00508379f $X=2.575 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A2_M1012_g N_A_165_74#_c_450_n 0.00109581f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A2_c_187_n N_A_264_74#_c_474_n 0.00124693f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A2_M1012_g N_A_264_74#_c_474_n 0.0151035f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A2_c_189_n N_A_264_74#_c_474_n 0.0247243f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A2_M1012_g N_A_264_74#_c_475_n 3.97481e-19 $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A2_M1012_g N_VGND_c_509_n 0.0124788f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A2_M1012_g N_VGND_c_515_n 0.00383152f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A2_M1012_g N_VGND_c_518_n 0.00757637f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A1_M1004_g N_A_27_368#_M1000_g 0.0233513f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_c_216_n N_A_27_368#_c_252_n 0.0382578f $X=3.145 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A1_M1004_g N_A_27_368#_c_252_n 9.38887e-19 $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A1_c_218_n N_A_27_368#_c_252_n 3.50433e-19 $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A1_c_216_n N_A_27_368#_c_296_n 0.0174338f $X=3.145 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A1_c_218_n N_A_27_368#_c_296_n 0.0250874f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A1_c_216_n N_A_27_368#_c_259_n 0.00365183f $X=3.145 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A1_c_218_n N_A_27_368#_c_259_n 0.00988402f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_183 N_A1_c_216_n N_A_27_368#_c_261_n 0.00170854f $X=3.145 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A1_M1004_g N_A_27_368#_c_261_n 5.96621e-19 $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A1_c_218_n N_A_27_368#_c_261_n 0.0231673f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A1_c_216_n N_VPWR_c_365_n 0.0174386f $X=3.145 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A1_c_216_n N_VPWR_c_369_n 0.0049405f $X=3.145 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A1_c_216_n N_VPWR_c_363_n 0.00508379f $X=3.145 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A1_c_216_n N_X_c_415_n 8.10615e-19 $X=3.145 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A1_c_216_n N_A_264_74#_c_474_n 3.13808e-19 $X=3.145 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A1_M1004_g N_A_264_74#_c_474_n 0.00351804f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_c_218_n N_A_264_74#_c_474_n 0.00993544f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_193 N_A1_M1004_g N_A_264_74#_c_475_n 0.00775604f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_M1004_g N_VGND_c_509_n 5.14838e-19 $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_c_216_n N_VGND_c_510_n 7.12986e-19 $X=3.145 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A1_M1004_g N_VGND_c_510_n 0.00657843f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A1_c_218_n N_VGND_c_510_n 0.00660905f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A1_M1004_g N_VGND_c_515_n 0.00434272f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A1_M1004_g N_VGND_c_518_n 0.0082141f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_27_368#_c_276_n N_VPWR_M1013_d 0.0257401f $X=2.065 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_201 N_A_27_368#_c_269_n N_VPWR_M1013_d 0.00666893f $X=0.775 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A_27_368#_c_296_n N_VPWR_M1009_d 0.0189236f $X=3.565 $Y=2.035 $X2=0
+ $Y2=0
cc_203 N_A_27_368#_c_259_n N_VPWR_M1009_d 0.00234639f $X=3.65 $Y=1.95 $X2=0
+ $Y2=0
cc_204 N_A_27_368#_c_265_n N_VPWR_c_364_n 0.0222698f $X=0.28 $Y=2.695 $X2=0
+ $Y2=0
cc_205 N_A_27_368#_c_267_n N_VPWR_c_364_n 0.0175483f $X=2.23 $Y=2.375 $X2=0
+ $Y2=0
cc_206 N_A_27_368#_c_269_n N_VPWR_c_364_n 0.067823f $X=0.775 $Y=1.97 $X2=0 $Y2=0
cc_207 N_A_27_368#_c_252_n N_VPWR_c_365_n 0.0105822f $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_27_368#_c_296_n N_VPWR_c_365_n 0.0258451f $X=3.565 $Y=2.035 $X2=0
+ $Y2=0
cc_209 N_A_27_368#_c_264_n N_VPWR_c_367_n 0.00954146f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_210 N_A_27_368#_c_265_n N_VPWR_c_368_n 0.0097982f $X=0.28 $Y=2.695 $X2=0
+ $Y2=0
cc_211 N_A_27_368#_c_267_n N_VPWR_c_369_n 0.0097982f $X=2.23 $Y=2.375 $X2=0
+ $Y2=0
cc_212 N_A_27_368#_c_252_n N_VPWR_c_370_n 0.00445602f $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A_27_368#_c_264_n N_VPWR_c_370_n 0.00411612f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A_27_368#_c_252_n N_VPWR_c_363_n 0.00861719f $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_A_27_368#_c_264_n N_VPWR_c_363_n 0.00751023f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_216 N_A_27_368#_c_265_n N_VPWR_c_363_n 0.0111907f $X=0.28 $Y=2.695 $X2=0
+ $Y2=0
cc_217 N_A_27_368#_c_267_n N_VPWR_c_363_n 0.0111907f $X=2.23 $Y=2.375 $X2=0
+ $Y2=0
cc_218 N_A_27_368#_c_276_n A_332_368# 0.00747797f $X=2.065 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_219 N_A_27_368#_c_296_n A_530_368# 0.0205616f $X=3.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_220 N_A_27_368#_c_252_n N_X_c_415_n 0.012608f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A_27_368#_c_264_n N_X_c_415_n 0.0130738f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A_27_368#_c_252_n N_X_c_416_n 0.00285426f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A_27_368#_c_253_n N_X_c_416_n 0.00277677f $X=4.095 $Y=1.395 $X2=0 $Y2=0
cc_224 N_A_27_368#_c_264_n N_X_c_416_n 0.00240464f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A_27_368#_c_259_n N_X_c_416_n 0.00565815f $X=3.65 $Y=1.95 $X2=0 $Y2=0
cc_226 N_A_27_368#_c_261_n N_X_c_416_n 0.00153915f $X=3.76 $Y=1.485 $X2=0 $Y2=0
cc_227 N_A_27_368#_M1000_g N_X_c_412_n 8.79499e-19 $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_27_368#_c_252_n N_X_c_412_n 0.00206544f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A_27_368#_M1007_g N_X_c_412_n 0.00708533f $X=4.17 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A_27_368#_c_255_n N_X_c_412_n 0.0100858f $X=4.295 $Y=1.675 $X2=0 $Y2=0
cc_231 N_A_27_368#_c_264_n N_X_c_412_n 0.00787412f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_27_368#_c_256_n N_X_c_412_n 0.0110677f $X=4.24 $Y=1.395 $X2=0 $Y2=0
cc_233 N_A_27_368#_c_259_n N_X_c_412_n 0.00535848f $X=3.65 $Y=1.95 $X2=0 $Y2=0
cc_234 N_A_27_368#_c_261_n N_X_c_412_n 0.0243803f $X=3.76 $Y=1.485 $X2=0 $Y2=0
cc_235 N_A_27_368#_M1000_g N_X_c_413_n 0.00675574f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_27_368#_M1007_g N_X_c_413_n 0.0177451f $X=4.17 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A_27_368#_M1000_g X 0.00303662f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_27_368#_c_252_n X 0.00426607f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_27_368#_M1007_g X 0.00692602f $X=4.17 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_27_368#_c_261_n X 0.0102861f $X=3.76 $Y=1.485 $X2=0 $Y2=0
cc_241 N_A_27_368#_c_257_n N_A_165_74#_c_449_n 0.0593848f $X=0.535 $Y=0.515
+ $X2=0 $Y2=0
cc_242 N_A_27_368#_M1000_g N_A_264_74#_c_474_n 2.49809e-19 $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_27_368#_c_258_n N_A_264_74#_c_476_n 0.00142925f $X=0.69 $Y=1.82 $X2=0
+ $Y2=0
cc_244 N_A_27_368#_M1000_g N_VGND_c_510_n 0.00805013f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_27_368#_c_252_n N_VGND_c_510_n 5.53507e-19 $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_246 N_A_27_368#_c_261_n N_VGND_c_510_n 0.00431466f $X=3.76 $Y=1.485 $X2=0
+ $Y2=0
cc_247 N_A_27_368#_M1007_g N_VGND_c_512_n 0.00925276f $X=4.17 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_27_368#_c_257_n N_VGND_c_513_n 0.0176636f $X=0.535 $Y=0.515 $X2=0
+ $Y2=0
cc_249 N_A_27_368#_M1000_g N_VGND_c_517_n 0.00434272f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A_27_368#_M1007_g N_VGND_c_517_n 0.00291513f $X=4.17 $Y=0.74 $X2=0
+ $Y2=0
cc_251 N_A_27_368#_M1000_g N_VGND_c_518_n 0.00821312f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_252 N_A_27_368#_M1007_g N_VGND_c_518_n 0.00363054f $X=4.17 $Y=0.74 $X2=0
+ $Y2=0
cc_253 N_A_27_368#_c_257_n N_VGND_c_518_n 0.0143978f $X=0.535 $Y=0.515 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_365_n N_X_c_415_n 0.027028f $X=3.57 $Y=2.455 $X2=0 $Y2=0
cc_255 N_VPWR_c_370_n N_X_c_415_n 0.0158009f $X=4.435 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_c_363_n N_X_c_415_n 0.0129424f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_367_n N_X_c_416_n 0.0887573f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_258 N_X_c_413_n N_VGND_c_510_n 0.0324855f $X=3.955 $Y=0.515 $X2=0 $Y2=0
cc_259 N_X_c_413_n N_VGND_c_512_n 0.0317393f $X=3.955 $Y=0.515 $X2=0 $Y2=0
cc_260 N_X_c_413_n N_VGND_c_517_n 0.0205856f $X=3.955 $Y=0.515 $X2=0 $Y2=0
cc_261 N_X_c_413_n N_VGND_c_518_n 0.0166302f $X=3.955 $Y=0.515 $X2=0 $Y2=0
cc_262 N_A_165_74#_c_448_n N_A_264_74#_M1010_d 0.00321664f $X=1.8 $Y=0.435
+ $X2=-0.19 $Y2=-0.245
cc_263 N_A_165_74#_M1003_d N_A_264_74#_c_474_n 0.0030579f $X=1.825 $Y=0.37 $X2=0
+ $Y2=0
cc_264 N_A_165_74#_c_448_n N_A_264_74#_c_474_n 0.00356375f $X=1.8 $Y=0.435 $X2=0
+ $Y2=0
cc_265 N_A_165_74#_c_450_n N_A_264_74#_c_474_n 0.020435f $X=1.965 $Y=0.435 $X2=0
+ $Y2=0
cc_266 N_A_165_74#_c_448_n N_A_264_74#_c_476_n 0.0127762f $X=1.8 $Y=0.435 $X2=0
+ $Y2=0
cc_267 N_A_165_74#_c_449_n N_A_264_74#_c_476_n 0.0124866f $X=1.03 $Y=0.515 $X2=0
+ $Y2=0
cc_268 N_A_165_74#_c_450_n N_VGND_c_509_n 0.0323609f $X=1.965 $Y=0.435 $X2=0
+ $Y2=0
cc_269 N_A_165_74#_c_448_n N_VGND_c_513_n 0.0269436f $X=1.8 $Y=0.435 $X2=0 $Y2=0
cc_270 N_A_165_74#_c_449_n N_VGND_c_513_n 0.00758556f $X=1.03 $Y=0.515 $X2=0
+ $Y2=0
cc_271 N_A_165_74#_c_450_n N_VGND_c_513_n 0.0142041f $X=1.965 $Y=0.435 $X2=0
+ $Y2=0
cc_272 N_A_165_74#_c_448_n N_VGND_c_518_n 0.0229064f $X=1.8 $Y=0.435 $X2=0 $Y2=0
cc_273 N_A_165_74#_c_449_n N_VGND_c_518_n 0.00627867f $X=1.03 $Y=0.515 $X2=0
+ $Y2=0
cc_274 N_A_165_74#_c_450_n N_VGND_c_518_n 0.011859f $X=1.965 $Y=0.435 $X2=0
+ $Y2=0
cc_275 N_A_264_74#_c_474_n N_VGND_M1012_s 0.0030579f $X=2.87 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A_264_74#_c_474_n N_VGND_c_509_n 0.02102f $X=2.87 $Y=1.095 $X2=0 $Y2=0
cc_277 N_A_264_74#_c_475_n N_VGND_c_509_n 0.0179318f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_278 N_A_264_74#_c_474_n N_VGND_c_510_n 0.00584871f $X=2.87 $Y=1.095 $X2=0
+ $Y2=0
cc_279 N_A_264_74#_c_475_n N_VGND_c_510_n 0.0244878f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_280 N_A_264_74#_c_475_n N_VGND_c_515_n 0.0109942f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_281 N_A_264_74#_c_475_n N_VGND_c_518_n 0.00904371f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
