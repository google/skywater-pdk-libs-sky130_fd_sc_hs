* File: sky130_fd_sc_hs__dfrbp_2.spice
* Created: Thu Aug 27 20:38:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfrbp_2.pex.spice"
.subckt sky130_fd_sc_hs__dfrbp_2  VNB VPB D RESET_B CLK VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1014 A_156_74# N_D_M1014_g N_A_70_74#_M1014_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1176 PD=0.66 PS=1.4 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_RESET_B_M1015_g A_156_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0821897 AS=0.0504 PD=0.78931 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_331_392#_M1003_d N_A_298_294#_M1003_g N_VGND_M1015_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.14481 PD=2.05 PS=1.39069 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1030 A_536_81# N_RESET_B_M1030_g N_VGND_M1030_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1281 PD=0.66 PS=1.45 NRD=18.564 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_614_81#_M1017_d N_A_331_392#_M1017_g A_536_81# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1281 AS=0.0504 PD=1.45 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_298_294#_M1004_d N_A_728_331#_M1004_g N_A_70_74#_M1004_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1456 PD=0.7 PS=1.63 NRD=0 NRS=25.704 M=1 R=2.8
+ SA=75000.3 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1035 N_A_614_81#_M1035_d N_A_818_418#_M1035_g N_A_298_294#_M1004_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.2184 AS=0.0588 PD=1.88 PS=0.7 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_A_728_331#_M1033_g N_A_818_418#_M1033_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.3983 AS=0.1998 PD=2.005 PS=2.02 NRD=78.36 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1005 N_A_728_331#_M1005_d N_CLK_M1005_g N_VGND_M1033_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.3983 PD=2.05 PS=2.005 NRD=0 NRS=78.36 M=1 R=4.93333
+ SA=75001.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_A_1586_149#_M1022_d N_A_728_331#_M1022_g N_A_1499_149#_M1022_s VNB
+ NLOWVT L=0.15 W=0.42 AD=0.0783879 AS=0.1197 PD=0.771207 PS=1.41 NRD=5.712
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1029 N_A_331_392#_M1029_d N_A_818_418#_M1029_g N_A_1586_149#_M1022_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.31255 AS=0.138112 PD=2.62 PS=1.35879 NRD=59.568
+ NRS=4.044 M=1 R=4.93333 SA=75000.5 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_1800_291#_M1010_g N_A_1499_149#_M1010_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1155 PD=0.7 PS=1.39 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1026 A_1974_74# N_RESET_B_M1026_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_A_1800_291#_M1023_d N_A_1586_149#_M1023_g A_1974_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_1586_149#_M1012_g N_Q_N_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1036 N_VGND_M1036_d N_A_1586_149#_M1036_g N_Q_N_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.124942 AS=0.1036 PD=1.14217 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1027 N_A_2363_352#_M1027_d N_A_1586_149#_M1027_g N_VGND_M1036_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1728 AS=0.108058 PD=1.82 PS=0.987826 NRD=0 NRS=7.488 M=1
+ R=4.26667 SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_Q_M1000_d N_A_2363_352#_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1019 N_Q_M1000_d N_A_2363_352#_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_70_74#_M1006_d N_D_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.1449 PD=0.72 PS=1.53 NRD=4.6886 NRS=28.1316 M=1 R=2.8 SA=75000.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_RESET_B_M1020_g N_A_70_74#_M1006_d VPB PSHORT L=0.15
+ W=0.42 AD=0.228175 AS=0.063 PD=1.59718 PS=0.72 NRD=229.013 NRS=4.6886 M=1
+ R=2.8 SA=75000.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_331_392#_M1001_d N_A_298_294#_M1001_g N_VPWR_M1020_d VPB PSHORT
+ L=0.15 W=1 AD=0.295 AS=0.543275 PD=2.59 PS=3.80282 NRD=1.9503 NRS=96.1754 M=1
+ R=6.66667 SA=75000.8 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1031 N_VPWR_M1031_d N_RESET_B_M1031_g N_A_298_294#_M1031_s VPB PSHORT L=0.15
+ W=0.42 AD=0.141475 AS=0.1176 PD=1.12 PS=1.4 NRD=114.91 NRS=4.6886 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1025 A_683_485# N_A_331_392#_M1025_g N_VPWR_M1031_d VPB PSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.141475 PD=0.66 PS=1.12 NRD=30.4759 NRS=46.886 M=1 R=2.8
+ SA=75001 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 N_A_298_294#_M1007_d N_A_728_331#_M1007_g A_683_485# VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.0504 PD=0.72 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75001.4 SB=75001 A=0.063 P=1.14 MULT=1
MM1013 N_A_70_74#_M1013_d N_A_818_418#_M1013_g N_A_298_294#_M1007_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.2793 AS=0.063 PD=2.17 PS=0.72 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75001.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_728_331#_M1008_g N_A_818_418#_M1008_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.372225 AS=0.3304 PD=1.805 PS=2.83 NRD=32.5247 NRS=1.7533
+ M=1 R=7.46667 SA=75000.2 SB=75001 A=0.168 P=2.54 MULT=1
MM1024 N_A_728_331#_M1024_d N_CLK_M1024_g N_VPWR_M1008_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.372225 PD=2.83 PS=1.805 NRD=1.7533 NRS=32.5247 M=1
+ R=7.46667 SA=75001 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1037 N_A_1586_149#_M1037_d N_A_728_331#_M1037_g N_A_331_392#_M1037_s VPB
+ PSHORT L=0.15 W=1 AD=0.265 AS=0.28 PD=2.15493 PS=2.56 NRD=47.2603 NRS=1.9503
+ M=1 R=6.66667 SA=75000.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1021 A_1755_389# N_A_818_418#_M1021_g N_A_1586_149#_M1037_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1113 PD=0.69 PS=0.90507 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.9 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1028 N_VPWR_M1028_d N_A_1800_291#_M1028_g A_1755_389# VPB PSHORT L=0.15 W=0.42
+ AD=0.1426 AS=0.0567 PD=1.155 PS=0.69 NRD=133.448 NRS=37.5088 M=1 R=2.8
+ SA=75001.3 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1016 N_A_1800_291#_M1016_d N_RESET_B_M1016_g N_VPWR_M1028_d VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.1426 PD=0.72 PS=1.155 NRD=4.6886 NRS=133.448 M=1 R=2.8
+ SA=75002 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_1586_149#_M1032_g N_A_1800_291#_M1016_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.0989045 AS=0.063 PD=0.820909 PS=0.72 NRD=46.886 NRS=4.6886
+ M=1 R=2.8 SA=75002.4 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1002 N_Q_N_M1002_d N_A_1586_149#_M1002_g N_VPWR_M1032_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.263745 PD=1.42 PS=2.18909 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.2 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1009 N_Q_N_M1002_d N_A_1586_149#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.222098 PD=1.42 PS=1.59019 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.7 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1034 N_A_2363_352#_M1034_d N_A_1586_149#_M1034_g N_VPWR_M1009_s VPB PSHORT
+ L=0.15 W=1 AD=0.39 AS=0.198302 PD=2.78 PS=1.41981 NRD=20.685 NRS=19.0302 M=1
+ R=6.66667 SA=75002.3 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1011 N_Q_M1011_d N_A_2363_352#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1018 N_Q_M1011_d N_A_2363_352#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75000.3 A=0.168 P=2.54 MULT=1
DX38_noxref VNB VPB NWDIODE A=25.4976 P=33.65
*
.include "sky130_fd_sc_hs__dfrbp_2.pxi.spice"
*
.ends
*
*
