* File: sky130_fd_sc_hs__a2bb2o_4.spice
* Created: Thu Aug 27 20:27:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a2bb2o_4.pex.spice"
.subckt sky130_fd_sc_hs__a2bb2o_4  VNB VPB A1_N A2_N B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_162_48#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_162_48#_M1007_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1007_d N_A_162_48#_M1010_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_162_48#_M1017_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=1.36203 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1012 N_A_586_94#_M1012_d N_A1_N_M1012_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.17797 NRD=0 NRS=46.872 M=1 R=4.26667
+ SA=75002.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_A2_N_M1020_g N_A_586_94#_M1012_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.309101 AS=0.0896 PD=1.61391 PS=0.92 NRD=53.436 NRS=0 M=1 R=4.26667
+ SA=75002.6 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1013 N_A_162_48#_M1013_d N_A_586_94#_M1013_g N_VGND_M1020_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.357399 PD=2.01 PS=1.86609 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_1009_74#_M1003_d N_B2_M1003_g N_A_162_48#_M1003_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1011 N_A_1009_74#_M1011_d N_B2_M1011_g N_A_162_48#_M1003_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_A_1009_74#_M1011_d N_B1_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=3.744 M=1 R=4.26667 SA=75001.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1008 N_A_1009_74#_M1008_d N_B1_M1008_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1024 PD=1.81 PS=0.96 NRD=0 NRS=3.744 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_162_48#_M1000_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_162_48#_M1015_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1015_d N_A_162_48#_M1018_g N_X_M1018_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1021_d N_A_162_48#_M1021_g N_X_M1018_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2184 AS=0.168 PD=1.51 PS=1.42 NRD=14.0658 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1004 A_583_368# N_A1_N_M1004_g N_VPWR_M1021_d VPB PSHORT L=0.15 W=1.12
+ AD=0.1344 AS=0.2184 PD=1.36 PS=1.51 NRD=11.426 NRS=5.2599 M=1 R=7.46667
+ SA=75002.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1001 N_A_586_94#_M1001_d N_A2_N_M1001_g A_583_368# VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.1344 PD=2.79 PS=1.36 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75002.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_A_162_48#_M1005_d N_A_586_94#_M1005_g N_A_820_392#_M1005_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1009 N_A_162_48#_M1005_d N_A_586_94#_M1009_g N_A_820_392#_M1009_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75002 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_B2_M1014_g N_A_820_392#_M1009_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1014_d N_B2_M1016_g N_A_820_392#_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_B1_M1019_g N_A_820_392#_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1019_d N_B1_M1022_g N_A_820_392#_M1022_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX23_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_hs__a2bb2o_4.pxi.spice"
*
.ends
*
*
