* File: sky130_fd_sc_hs__a22o_2.pxi.spice
* Created: Tue Sep  1 19:51:12 2020
* 
x_PM_SKY130_FD_SC_HS__A22O_2%A_81_48# N_A_81_48#_M1009_d N_A_81_48#_M1004_d
+ N_A_81_48#_c_66_n N_A_81_48#_M1000_g N_A_81_48#_c_73_n N_A_81_48#_M1001_g
+ N_A_81_48#_c_67_n N_A_81_48#_M1010_g N_A_81_48#_c_74_n N_A_81_48#_M1002_g
+ N_A_81_48#_c_75_n N_A_81_48#_c_68_n N_A_81_48#_c_69_n N_A_81_48#_c_80_p
+ N_A_81_48#_c_104_p N_A_81_48#_c_94_p N_A_81_48#_c_70_n N_A_81_48#_c_71_n
+ N_A_81_48#_c_72_n N_A_81_48#_c_92_p PM_SKY130_FD_SC_HS__A22O_2%A_81_48#
x_PM_SKY130_FD_SC_HS__A22O_2%A1 N_A1_c_144_n N_A1_M1003_g N_A1_M1009_g A1
+ N_A1_c_146_n PM_SKY130_FD_SC_HS__A22O_2%A1
x_PM_SKY130_FD_SC_HS__A22O_2%B1 N_B1_c_178_n N_B1_M1004_g N_B1_M1007_g B1
+ N_B1_c_180_n PM_SKY130_FD_SC_HS__A22O_2%B1
x_PM_SKY130_FD_SC_HS__A22O_2%B2 N_B2_M1011_g N_B2_c_212_n N_B2_M1005_g B2
+ PM_SKY130_FD_SC_HS__A22O_2%B2
x_PM_SKY130_FD_SC_HS__A22O_2%A2 N_A2_M1006_g N_A2_c_241_n N_A2_M1008_g A2
+ N_A2_c_242_n PM_SKY130_FD_SC_HS__A22O_2%A2
x_PM_SKY130_FD_SC_HS__A22O_2%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1008_d
+ N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n
+ N_VPWR_c_269_n VPWR N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n
+ N_VPWR_c_263_n PM_SKY130_FD_SC_HS__A22O_2%VPWR
x_PM_SKY130_FD_SC_HS__A22O_2%X N_X_M1000_s N_X_M1001_d N_X_c_313_n N_X_c_310_n
+ N_X_c_316_n X X X X X N_X_c_312_n PM_SKY130_FD_SC_HS__A22O_2%X
x_PM_SKY130_FD_SC_HS__A22O_2%A_388_368# N_A_388_368#_M1003_d
+ N_A_388_368#_M1005_d N_A_388_368#_c_342_n N_A_388_368#_c_338_n
+ N_A_388_368#_c_339_n N_A_388_368#_c_340_n
+ PM_SKY130_FD_SC_HS__A22O_2%A_388_368#
x_PM_SKY130_FD_SC_HS__A22O_2%VGND N_VGND_M1000_d N_VGND_M1010_d N_VGND_M1011_d
+ N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n N_VGND_c_370_n
+ N_VGND_c_371_n VGND N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n
+ N_VGND_c_375_n PM_SKY130_FD_SC_HS__A22O_2%VGND
x_PM_SKY130_FD_SC_HS__A22O_2%A_304_74# N_A_304_74#_M1009_s N_A_304_74#_M1006_d
+ N_A_304_74#_c_412_n N_A_304_74#_c_413_n N_A_304_74#_c_414_n
+ N_A_304_74#_c_451_p N_A_304_74#_c_415_n N_A_304_74#_c_416_n
+ N_A_304_74#_c_417_n PM_SKY130_FD_SC_HS__A22O_2%A_304_74#
cc_1 VNB N_A_81_48#_c_66_n 0.0199307f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.22
cc_2 VNB N_A_81_48#_c_67_n 0.0176642f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.22
cc_3 VNB N_A_81_48#_c_68_n 0.0167228f $X=-0.19 $Y=-0.245 $X2=2 $Y2=1.095
cc_4 VNB N_A_81_48#_c_69_n 0.00613798f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.095
cc_5 VNB N_A_81_48#_c_70_n 7.42537e-19 $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.385
cc_6 VNB N_A_81_48#_c_71_n 0.10555f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.385
cc_7 VNB N_A_81_48#_c_72_n 0.00233643f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.55
cc_8 VNB N_A1_c_144_n 0.0242699f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=0.37
cc_9 VNB N_A1_M1009_g 0.0275155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_146_n 0.00392334f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_11 VNB N_B1_c_178_n 0.0227068f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=0.37
cc_12 VNB N_B1_M1007_g 0.0237683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_180_n 0.00472951f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_14 VNB N_B2_M1011_g 0.0251119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_c_212_n 0.0215738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB B2 0.00585622f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_17 VNB N_A2_M1006_g 0.0345407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_241_n 0.0473054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_242_n 0.00404344f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_20 VNB N_VPWR_c_263_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB X 0.00650146f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_22 VNB N_VGND_c_366_n 0.0101995f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.765
cc_23 VNB N_VGND_c_367_n 0.0511447f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_24 VNB N_VGND_c_368_n 0.0134317f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.765
cc_25 VNB N_VGND_c_369_n 0.00941023f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.385
cc_26 VNB N_VGND_c_370_n 0.0389074f $X=-0.19 $Y=-0.245 $X2=2 $Y2=1.095
cc_27 VNB N_VGND_c_371_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.095
cc_28 VNB N_VGND_c_372_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=2.165 $Y2=1.01
cc_29 VNB N_VGND_c_373_n 0.0199471f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.492
cc_30 VNB N_VGND_c_374_n 0.237175f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.492
cc_31 VNB N_VGND_c_375_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_304_74#_c_412_n 0.00370491f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_33 VNB N_A_304_74#_c_413_n 0.0048983f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_34 VNB N_A_304_74#_c_414_n 0.00412286f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_35 VNB N_A_304_74#_c_415_n 0.0137f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_36 VNB N_A_304_74#_c_416_n 0.00735846f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.765
cc_37 VNB N_A_304_74#_c_417_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.18
cc_38 VPB N_A_81_48#_c_73_n 0.0165358f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=1.765
cc_39 VPB N_A_81_48#_c_74_n 0.0164337f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=1.765
cc_40 VPB N_A_81_48#_c_75_n 0.00124183f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=1.95
cc_41 VPB N_A_81_48#_c_71_n 0.0143663f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.385
cc_42 VPB N_A1_c_144_n 0.0262143f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=0.37
cc_43 VPB N_A1_c_146_n 0.00263019f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_44 VPB N_B1_c_178_n 0.0249146f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=0.37
cc_45 VPB N_B1_c_180_n 0.00402621f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_46 VPB N_B2_c_212_n 0.0256491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB B2 0.006451f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=0.74
cc_48 VPB N_A2_c_241_n 0.0372068f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A2_c_242_n 0.00703186f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_50 VPB N_VPWR_c_264_n 0.0458691f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_51 VPB N_VPWR_c_265_n 0.00731821f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=1.765
cc_52 VPB N_VPWR_c_266_n 0.0121909f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=2.4
cc_53 VPB N_VPWR_c_267_n 0.0519518f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.385
cc_54 VPB N_VPWR_c_268_n 0.017577f $X=-0.19 $Y=1.66 $X2=2 $Y2=1.095
cc_55 VPB N_VPWR_c_269_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.415 $Y2=1.095
cc_56 VPB N_VPWR_c_270_n 0.0182909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_271_n 0.0411787f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.385
cc_58 VPB N_VPWR_c_272_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=1.492
cc_59 VPB N_VPWR_c_263_n 0.0876923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_X_c_310_n 0.00217048f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_61 VPB X 0.00296132f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=0.74
cc_62 VPB N_X_c_312_n 0.00952671f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.115
cc_63 VPB N_A_388_368#_c_338_n 0.0150135f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_64 VPB N_A_388_368#_c_339_n 0.00323592f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_65 VPB N_A_388_368#_c_340_n 7.13292e-19 $X=-0.19 $Y=1.66 $X2=0.91 $Y2=0.74
cc_66 N_A_81_48#_c_74_n N_A1_c_144_n 0.0223501f $X=1.325 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_67 N_A_81_48#_c_75_n N_A1_c_144_n 0.00145794f $X=1.33 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_68 N_A_81_48#_c_68_n N_A1_c_144_n 0.00126708f $X=2 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_69 N_A_81_48#_c_80_p N_A1_c_144_n 0.0170704f $X=2.455 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_70 N_A_81_48#_c_70_n N_A1_c_144_n 3.80775e-19 $X=1.25 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_81_48#_c_71_n N_A1_c_144_n 0.0235088f $X=1.25 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_81_48#_c_68_n N_A1_M1009_g 0.0160323f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_73 N_A_81_48#_c_70_n N_A1_M1009_g 0.0019081f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_74 N_A_81_48#_c_71_n N_A1_M1009_g 0.00473768f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_75 N_A_81_48#_c_68_n N_A1_c_146_n 0.0243073f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_76 N_A_81_48#_c_80_p N_A1_c_146_n 0.0226059f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_77 N_A_81_48#_c_70_n N_A1_c_146_n 0.0330964f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_78 N_A_81_48#_c_71_n N_A1_c_146_n 0.00250676f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_79 N_A_81_48#_c_68_n N_B1_c_178_n 0.00351433f $X=2 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_81_48#_c_80_p N_B1_c_178_n 0.013077f $X=2.455 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_81 N_A_81_48#_c_92_p N_B1_c_178_n 0.00569691f $X=2.54 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_82 N_A_81_48#_c_68_n N_B1_M1007_g 0.00442568f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_81_48#_c_94_p N_B1_M1007_g 0.00514063f $X=2.165 $Y=0.76 $X2=0 $Y2=0
cc_84 N_A_81_48#_c_68_n N_B1_c_180_n 0.0219116f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_85 N_A_81_48#_c_80_p N_B1_c_180_n 0.025054f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_86 N_A_81_48#_c_92_p N_B1_c_180_n 0.00353587f $X=2.54 $Y=2.115 $X2=0 $Y2=0
cc_87 N_A_81_48#_c_80_p N_VPWR_M1002_s 0.010009f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A_81_48#_c_73_n N_VPWR_c_264_n 0.00998224f $X=0.875 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_81_48#_c_71_n N_VPWR_c_264_n 0.00150952f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_90 N_A_81_48#_c_73_n N_VPWR_c_265_n 5.55114e-19 $X=0.875 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_81_48#_c_74_n N_VPWR_c_265_n 0.012746f $X=1.325 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_81_48#_c_80_p N_VPWR_c_265_n 0.0209091f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_81_48#_c_104_p N_VPWR_c_265_n 0.00114279f $X=1.415 $Y=2.035 $X2=0
+ $Y2=0
cc_94 N_A_81_48#_c_73_n N_VPWR_c_270_n 0.00411612f $X=0.875 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_81_48#_c_74_n N_VPWR_c_270_n 0.00413917f $X=1.325 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_81_48#_c_73_n N_VPWR_c_263_n 0.00752331f $X=0.875 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A_81_48#_c_74_n N_VPWR_c_263_n 0.00817726f $X=1.325 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_81_48#_c_73_n N_X_c_313_n 0.00168175f $X=0.875 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_81_48#_c_74_n N_X_c_313_n 0.0025256f $X=1.325 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_81_48#_c_73_n N_X_c_310_n 0.0072148f $X=0.875 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A_81_48#_c_73_n N_X_c_316_n 0.0127177f $X=0.875 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_81_48#_c_74_n N_X_c_316_n 0.004142f $X=1.325 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A_81_48#_c_66_n X 0.0148558f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_104 N_A_81_48#_c_67_n X 0.0177235f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_105 N_A_81_48#_c_75_n X 0.00627104f $X=1.33 $Y=1.95 $X2=0 $Y2=0
cc_106 N_A_81_48#_c_69_n X 0.011439f $X=1.415 $Y=1.095 $X2=0 $Y2=0
cc_107 N_A_81_48#_c_70_n X 0.0222666f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_108 N_A_81_48#_c_71_n X 0.0434158f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_109 N_A_81_48#_c_73_n N_X_c_312_n 0.00987153f $X=0.875 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_81_48#_c_74_n N_X_c_312_n 4.77242e-19 $X=1.325 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_81_48#_c_75_n N_X_c_312_n 0.0117914f $X=1.33 $Y=1.95 $X2=0 $Y2=0
cc_112 N_A_81_48#_c_71_n N_X_c_312_n 0.00955127f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_113 N_A_81_48#_c_80_p N_A_388_368#_M1003_d 0.00606883f $X=2.455 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_114 N_A_81_48#_c_80_p N_A_388_368#_c_342_n 0.0171814f $X=2.455 $Y=2.035 $X2=0
+ $Y2=0
cc_115 N_A_81_48#_c_92_p N_A_388_368#_c_342_n 0.0298377f $X=2.54 $Y=2.115 $X2=0
+ $Y2=0
cc_116 N_A_81_48#_c_92_p N_A_388_368#_c_338_n 0.0183738f $X=2.54 $Y=2.115 $X2=0
+ $Y2=0
cc_117 N_A_81_48#_c_74_n N_A_388_368#_c_339_n 4.80813e-19 $X=1.325 $Y=1.765
+ $X2=0 $Y2=0
cc_118 N_A_81_48#_c_69_n N_VGND_M1010_d 0.0030302f $X=1.415 $Y=1.095 $X2=0 $Y2=0
cc_119 N_A_81_48#_c_66_n N_VGND_c_367_n 0.00647412f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_120 N_A_81_48#_c_67_n N_VGND_c_368_n 0.00698798f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_121 N_A_81_48#_c_69_n N_VGND_c_368_n 0.0182898f $X=1.415 $Y=1.095 $X2=0 $Y2=0
cc_122 N_A_81_48#_c_71_n N_VGND_c_368_n 0.00259377f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_123 N_A_81_48#_c_66_n N_VGND_c_372_n 0.00434272f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_124 N_A_81_48#_c_67_n N_VGND_c_372_n 0.00434272f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_125 N_A_81_48#_c_66_n N_VGND_c_374_n 0.00823889f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_126 N_A_81_48#_c_67_n N_VGND_c_374_n 0.00825283f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_127 N_A_81_48#_c_68_n N_A_304_74#_M1009_s 0.00271234f $X=2 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_81_48#_c_68_n N_A_304_74#_c_412_n 0.021673f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_129 N_A_81_48#_M1009_d N_A_304_74#_c_413_n 0.00250873f $X=1.955 $Y=0.37 $X2=0
+ $Y2=0
cc_130 N_A_81_48#_c_68_n N_A_304_74#_c_413_n 0.00304353f $X=2 $Y=1.095 $X2=0
+ $Y2=0
cc_131 N_A_81_48#_c_94_p N_A_304_74#_c_413_n 0.0194097f $X=2.165 $Y=0.76 $X2=0
+ $Y2=0
cc_132 N_A_81_48#_c_68_n N_A_304_74#_c_416_n 0.0104256f $X=2 $Y=1.095 $X2=0
+ $Y2=0
cc_133 N_A1_c_144_n N_B1_c_178_n 0.0477579f $X=1.865 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A1_c_146_n N_B1_c_178_n 4.06432e-19 $X=1.79 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A1_M1009_g N_B1_M1007_g 0.0301069f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A1_c_144_n N_B1_c_180_n 0.00276327f $X=1.865 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A1_c_146_n N_B1_c_180_n 0.034584f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A1_c_144_n N_VPWR_c_265_n 0.00621193f $X=1.865 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A1_c_144_n N_VPWR_c_271_n 0.00451897f $X=1.865 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A1_c_144_n N_VPWR_c_263_n 0.00457541f $X=1.865 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_144_n N_A_388_368#_c_342_n 0.00744575f $X=1.865 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A1_c_144_n N_A_388_368#_c_339_n 0.00174271f $X=1.865 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A1_M1009_g N_VGND_c_368_n 0.00174891f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_M1009_g N_VGND_c_370_n 0.00278247f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A1_M1009_g N_VGND_c_374_n 0.00359137f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A1_M1009_g N_A_304_74#_c_412_n 0.00730569f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A1_M1009_g N_A_304_74#_c_413_n 0.008259f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A1_M1009_g N_A_304_74#_c_414_n 0.00395315f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_149 N_B1_M1007_g N_B2_M1011_g 0.0500418f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_150 N_B1_c_178_n N_B2_c_212_n 0.0492579f $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_151 N_B1_c_180_n N_B2_c_212_n 7.86793e-19 $X=2.33 $Y=1.515 $X2=0 $Y2=0
cc_152 N_B1_c_178_n B2 7.46006e-19 $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_153 N_B1_c_180_n B2 0.0297654f $X=2.33 $Y=1.515 $X2=0 $Y2=0
cc_154 N_B1_c_178_n N_VPWR_c_271_n 7.44201e-19 $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_155 N_B1_c_178_n N_A_388_368#_c_342_n 0.00866602f $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_B1_c_178_n N_A_388_368#_c_338_n 0.00981448f $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_157 N_B1_c_178_n N_A_388_368#_c_339_n 0.00114023f $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_158 N_B1_c_178_n N_A_388_368#_c_340_n 5.87231e-19 $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_B1_M1007_g N_VGND_c_370_n 0.00278271f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_160 N_B1_M1007_g N_VGND_c_374_n 0.00353949f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_161 N_B1_M1007_g N_A_304_74#_c_412_n 4.62714e-19 $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_162 N_B1_M1007_g N_A_304_74#_c_413_n 0.0127288f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_163 N_B1_M1007_g N_A_304_74#_c_416_n 9.3266e-19 $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_164 N_B2_M1011_g N_A2_M1006_g 0.024575f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_165 N_B2_c_212_n N_A2_c_241_n 0.0422813f $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_166 B2 N_A2_c_241_n 0.0038009f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_167 N_B2_c_212_n N_A2_c_242_n 2.88866e-19 $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_168 B2 N_A2_c_242_n 0.035317f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_169 N_B2_c_212_n N_VPWR_c_267_n 2.84074e-19 $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_170 N_B2_c_212_n N_VPWR_c_271_n 7.44201e-19 $X=2.815 $Y=1.765 $X2=0 $Y2=0
cc_171 N_B2_c_212_n N_A_388_368#_c_342_n 6.34207e-19 $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_B2_c_212_n N_A_388_368#_c_338_n 0.0109883f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_173 N_B2_c_212_n N_A_388_368#_c_340_n 0.0122989f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_174 B2 N_A_388_368#_c_340_n 0.0271212f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_175 N_B2_M1011_g N_VGND_c_369_n 0.00225437f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B2_M1011_g N_VGND_c_370_n 0.00461464f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B2_M1011_g N_VGND_c_374_n 0.00908275f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_178 N_B2_M1011_g N_A_304_74#_c_413_n 0.00120883f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B2_M1011_g N_A_304_74#_c_415_n 0.014921f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B2_c_212_n N_A_304_74#_c_415_n 0.00418988f $X=2.815 $Y=1.765 $X2=0
+ $Y2=0
cc_181 B2 N_A_304_74#_c_415_n 0.0409488f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_182 N_B2_M1011_g N_A_304_74#_c_417_n 8.17877e-19 $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A2_c_241_n N_VPWR_c_267_n 0.0188061f $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A2_c_242_n N_VPWR_c_267_n 0.0256701f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A2_c_241_n N_VPWR_c_271_n 0.00443511f $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A2_c_241_n N_VPWR_c_263_n 0.00460931f $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A2_c_241_n N_A_388_368#_c_338_n 6.25105e-19 $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A2_c_241_n N_A_388_368#_c_340_n 0.00554206f $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A2_M1006_g N_VGND_c_369_n 0.00600897f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A2_M1006_g N_VGND_c_373_n 0.00434272f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A2_M1006_g N_VGND_c_374_n 0.00824829f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A2_M1006_g N_A_304_74#_c_415_n 0.018512f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A2_c_241_n N_A_304_74#_c_415_n 0.00285838f $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_A2_c_242_n N_A_304_74#_c_415_n 0.0253731f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A2_M1006_g N_A_304_74#_c_417_n 0.0102372f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_196 N_VPWR_c_265_n N_X_c_313_n 0.0466627f $X=1.55 $Y=2.375 $X2=0 $Y2=0
cc_197 N_VPWR_c_270_n N_X_c_310_n 0.0122783f $X=1.385 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_c_263_n N_X_c_310_n 0.0100573f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_264_n N_X_c_316_n 0.068395f $X=0.65 $Y=2.225 $X2=0 $Y2=0
cc_200 N_VPWR_M1001_s N_X_c_312_n 0.00486797f $X=0.525 $Y=1.84 $X2=0 $Y2=0
cc_201 N_VPWR_c_264_n N_X_c_312_n 0.0165971f $X=0.65 $Y=2.225 $X2=0 $Y2=0
cc_202 N_VPWR_c_265_n N_A_388_368#_c_342_n 0.0406488f $X=1.55 $Y=2.375 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_267_n N_A_388_368#_c_338_n 0.0147692f $X=3.56 $Y=2.115 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_271_n N_A_388_368#_c_338_n 0.0649714f $X=3.395 $Y=3.33 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_263_n N_A_388_368#_c_338_n 0.0369098f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_265_n N_A_388_368#_c_339_n 0.0126524f $X=1.55 $Y=2.375 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_271_n N_A_388_368#_c_339_n 0.0236566f $X=3.395 $Y=3.33 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_263_n N_A_388_368#_c_339_n 0.0128296f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_209 N_VPWR_c_267_n N_A_388_368#_c_340_n 0.0384784f $X=3.56 $Y=2.115 $X2=0
+ $Y2=0
cc_210 X N_VGND_c_367_n 0.0294122f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_211 X N_VGND_c_368_n 0.0182902f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_212 X N_VGND_c_372_n 0.0144922f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_213 X N_VGND_c_374_n 0.0118826f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_214 N_VGND_c_368_n N_A_304_74#_c_412_n 0.0291511f $X=1.125 $Y=0.675 $X2=0
+ $Y2=0
cc_215 N_VGND_c_369_n N_A_304_74#_c_413_n 0.00898192f $X=3.035 $Y=0.675 $X2=0
+ $Y2=0
cc_216 N_VGND_c_370_n N_A_304_74#_c_413_n 0.0544911f $X=2.87 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_374_n N_A_304_74#_c_413_n 0.0305408f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_368_n N_A_304_74#_c_414_n 0.0127054f $X=1.125 $Y=0.675 $X2=0
+ $Y2=0
cc_219 N_VGND_c_370_n N_A_304_74#_c_414_n 0.0233048f $X=2.87 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_374_n N_A_304_74#_c_414_n 0.0126653f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_M1011_d N_A_304_74#_c_415_n 0.00309832f $X=2.855 $Y=0.37 $X2=0
+ $Y2=0
cc_222 N_VGND_c_369_n N_A_304_74#_c_415_n 0.022455f $X=3.035 $Y=0.675 $X2=0
+ $Y2=0
cc_223 N_VGND_c_369_n N_A_304_74#_c_417_n 0.0191765f $X=3.035 $Y=0.675 $X2=0
+ $Y2=0
cc_224 N_VGND_c_373_n N_A_304_74#_c_417_n 0.0145639f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_374_n N_A_304_74#_c_417_n 0.0119984f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_226 N_A_304_74#_c_451_p A_491_74# 0.00196494f $X=2.585 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
