* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_1474_446# a_2320_410# VPB pshort w=840000u l=150000u
+  ad=2.9038e+12p pd=2.241e+07u as=2.31e+11p ps=2.23e+06u
M1001 Q_N a_1474_446# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.83492e+12p ps=1.558e+07u
M1002 a_1017_379# a_520_87# a_671_93# VPB pshort w=840000u l=150000u
+  ad=2.268e+11p pd=2.22e+06u as=3.276e+11p ps=2.46e+06u
M1003 a_520_87# a_27_74# a_422_125# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.7605e+11p ps=1.9e+06u
M1004 Q a_2320_410# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1005 a_1318_119# a_671_93# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1006 VGND RESET_B a_1062_93# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1007 a_713_379# a_27_74# a_520_87# VPB pshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.289e+11p ps=2.42e+06u
M1008 VPWR RESET_B a_1062_93# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1009 a_1474_446# SET_B VPWR VPB pshort w=1e+06u l=150000u
+  ad=3.65e+11p pd=2.73e+06u as=0p ps=0u
M1010 a_1311_424# a_214_74# a_1318_119# VNB nlowvt w=550000u l=150000u
+  ad=2.317e+11p pd=2.33e+06u as=0p ps=0u
M1011 a_1418_508# a_214_74# a_1311_424# VPB pshort w=420000u l=150000u
+  ad=1.239e+11p pd=1.43e+06u as=2.856e+11p ps=2.45e+06u
M1012 a_1498_74# a_27_74# a_1311_424# VNB nlowvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1013 a_214_74# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_1203_379# a_671_93# VPWR VPB pshort w=840000u l=150000u
+  ad=3.591e+11p pd=2.91e+06u as=0p ps=0u
M1015 a_214_74# a_27_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1016 VGND a_1474_446# a_2320_410# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1017 a_1814_392# a_1311_424# a_1474_446# VPB pshort w=1e+06u l=150000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1018 a_422_125# D VPWR VPB pshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1019 VGND a_1474_446# a_1498_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1474_446# a_1418_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_671_93# a_520_87# a_872_119# VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=6.465e+11p ps=4.96e+06u
M1022 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1023 a_520_87# a_214_74# a_422_125# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_606_87# a_214_74# a_520_87# VNB nlowvt w=420000u l=150000u
+  ad=1.645e+11p pd=1.81e+06u as=0p ps=0u
M1025 a_671_93# SET_B VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1311_424# a_27_74# a_1203_379# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1474_446# a_1311_424# a_1708_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=4.884e+11p ps=4.28e+06u
M1028 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1029 VPWR a_671_93# a_713_379# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_872_119# a_1062_93# a_671_93# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Q_N a_1474_446# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1032 a_1708_74# a_1062_93# a_1474_446# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_422_125# D VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_872_119# SET_B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1708_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_1062_93# a_1017_379# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_671_93# a_606_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Q a_2320_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1039 VPWR a_1062_93# a_1814_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
