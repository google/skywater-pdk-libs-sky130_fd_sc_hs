* File: sky130_fd_sc_hs__o2111ai_2.pxi.spice
* Created: Tue Sep  1 20:13:23 2020
* 
x_PM_SKY130_FD_SC_HS__O2111AI_2%D1 N_D1_c_105_n N_D1_M1018_g N_D1_c_100_n
+ N_D1_M1012_g N_D1_c_101_n N_D1_M1014_g N_D1_c_106_n N_D1_M1019_g N_D1_c_102_n
+ N_D1_c_103_n D1 PM_SKY130_FD_SC_HS__O2111AI_2%D1
x_PM_SKY130_FD_SC_HS__O2111AI_2%C1 N_C1_M1004_g N_C1_c_152_n N_C1_M1000_g
+ N_C1_M1005_g N_C1_c_153_n N_C1_M1016_g C1 N_C1_c_151_n
+ PM_SKY130_FD_SC_HS__O2111AI_2%C1
x_PM_SKY130_FD_SC_HS__O2111AI_2%B1 N_B1_c_214_n N_B1_M1002_g N_B1_c_207_n
+ N_B1_c_216_n N_B1_M1003_g N_B1_M1007_g N_B1_M1009_g N_B1_c_210_n N_B1_c_211_n
+ N_B1_c_212_n B1 B1 B1 PM_SKY130_FD_SC_HS__O2111AI_2%B1
x_PM_SKY130_FD_SC_HS__O2111AI_2%A2 N_A2_M1001_g N_A2_c_275_n N_A2_M1008_g
+ N_A2_M1015_g N_A2_c_276_n N_A2_M1011_g A2 A2 N_A2_c_274_n
+ PM_SKY130_FD_SC_HS__O2111AI_2%A2
x_PM_SKY130_FD_SC_HS__O2111AI_2%A1 N_A1_M1006_g N_A1_c_323_n N_A1_M1013_g
+ N_A1_M1010_g N_A1_c_324_n N_A1_M1017_g A1 A1 N_A1_c_322_n
+ PM_SKY130_FD_SC_HS__O2111AI_2%A1
x_PM_SKY130_FD_SC_HS__O2111AI_2%VPWR N_VPWR_M1018_s N_VPWR_M1019_s
+ N_VPWR_M1016_d N_VPWR_M1003_s N_VPWR_M1013_d N_VPWR_c_364_n N_VPWR_c_365_n
+ N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n
+ VPWR N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n
+ N_VPWR_c_363_n N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n
+ PM_SKY130_FD_SC_HS__O2111AI_2%VPWR
x_PM_SKY130_FD_SC_HS__O2111AI_2%Y N_Y_M1012_s N_Y_M1018_d N_Y_M1000_s
+ N_Y_M1002_d N_Y_M1008_d N_Y_c_450_n N_Y_c_444_n N_Y_c_445_n N_Y_c_471_n
+ N_Y_c_446_n N_Y_c_447_n N_Y_c_448_n N_Y_c_490_n N_Y_c_495_n Y Y Y Y Y
+ N_Y_c_443_n Y Y PM_SKY130_FD_SC_HS__O2111AI_2%Y
x_PM_SKY130_FD_SC_HS__O2111AI_2%A_697_368# N_A_697_368#_M1008_s
+ N_A_697_368#_M1011_s N_A_697_368#_M1017_s N_A_697_368#_c_529_n
+ N_A_697_368#_c_530_n N_A_697_368#_c_531_n N_A_697_368#_c_536_n
+ N_A_697_368#_c_555_n N_A_697_368#_c_537_n N_A_697_368#_c_532_n
+ N_A_697_368#_c_533_n PM_SKY130_FD_SC_HS__O2111AI_2%A_697_368#
x_PM_SKY130_FD_SC_HS__O2111AI_2%A_40_74# N_A_40_74#_M1012_d N_A_40_74#_M1014_d
+ N_A_40_74#_M1005_d N_A_40_74#_c_568_n N_A_40_74#_c_569_n N_A_40_74#_c_570_n
+ N_A_40_74#_c_571_n N_A_40_74#_c_572_n N_A_40_74#_c_586_n
+ PM_SKY130_FD_SC_HS__O2111AI_2%A_40_74#
x_PM_SKY130_FD_SC_HS__O2111AI_2%A_299_74# N_A_299_74#_M1004_s
+ N_A_299_74#_M1007_s N_A_299_74#_c_608_n N_A_299_74#_c_615_n
+ N_A_299_74#_c_609_n PM_SKY130_FD_SC_HS__O2111AI_2%A_299_74#
x_PM_SKY130_FD_SC_HS__O2111AI_2%A_510_74# N_A_510_74#_M1007_d
+ N_A_510_74#_M1009_d N_A_510_74#_M1015_d N_A_510_74#_M1010_d
+ N_A_510_74#_c_634_n N_A_510_74#_c_635_n N_A_510_74#_c_636_n
+ N_A_510_74#_c_637_n N_A_510_74#_c_638_n N_A_510_74#_c_639_n
+ N_A_510_74#_c_640_n N_A_510_74#_c_641_n N_A_510_74#_c_642_n
+ N_A_510_74#_c_643_n PM_SKY130_FD_SC_HS__O2111AI_2%A_510_74#
x_PM_SKY130_FD_SC_HS__O2111AI_2%VGND N_VGND_M1001_s N_VGND_M1006_s
+ N_VGND_c_697_n N_VGND_c_698_n VGND N_VGND_c_699_n N_VGND_c_700_n
+ N_VGND_c_701_n N_VGND_c_702_n N_VGND_c_703_n N_VGND_c_704_n
+ PM_SKY130_FD_SC_HS__O2111AI_2%VGND
cc_1 VNB N_D1_c_100_n 0.0204008f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.22
cc_2 VNB N_D1_c_101_n 0.0159551f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.22
cc_3 VNB N_D1_c_102_n 0.0507325f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_4 VNB N_D1_c_103_n 0.0500731f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.492
cc_5 VNB D1 0.0126727f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_C1_M1004_g 0.0219968f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_7 VNB N_C1_M1005_g 0.0275487f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_8 VNB C1 0.0105601f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.492
cc_9 VNB N_C1_c_151_n 0.0576224f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_10 VNB N_B1_c_207_n 0.0120923f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.22
cc_11 VNB N_B1_M1007_g 0.0314339f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_12 VNB N_B1_M1009_g 0.024203f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.492
cc_13 VNB N_B1_c_210_n 0.0147919f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.492
cc_14 VNB N_B1_c_211_n 0.0142678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_212_n 0.024603f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_16 VNB B1 0.00931452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_M1001_g 0.0232975f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_18 VNB N_A2_M1015_g 0.0232975f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_19 VNB A2 0.00232957f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.492
cc_20 VNB N_A2_c_274_n 0.0343051f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_21 VNB N_A1_M1006_g 0.0245199f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_22 VNB N_A1_M1010_g 0.0328675f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_23 VNB A1 0.0161791f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.492
cc_24 VNB N_A1_c_322_n 0.0453025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_363_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_443_n 0.00289639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_40_74#_c_568_n 0.0222939f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_28 VNB N_A_40_74#_c_569_n 0.00448726f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.492
cc_29 VNB N_A_40_74#_c_570_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.492
cc_30 VNB N_A_40_74#_c_571_n 0.00325f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.492
cc_31 VNB N_A_40_74#_c_572_n 0.0157968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_299_74#_c_608_n 0.0199129f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.22
cc_33 VNB N_A_299_74#_c_609_n 0.00240543f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_34 VNB N_A_510_74#_c_634_n 0.00380647f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.492
cc_35 VNB N_A_510_74#_c_635_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.492
cc_36 VNB N_A_510_74#_c_636_n 0.00417749f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_37 VNB N_A_510_74#_c_637_n 0.00178889f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_38 VNB N_A_510_74#_c_638_n 0.00575126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_510_74#_c_639_n 0.00207041f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_40 VNB N_A_510_74#_c_640_n 0.0148256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_510_74#_c_641_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_510_74#_c_642_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_510_74#_c_643_n 0.00211286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_697_n 0.00335558f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.74
cc_45 VNB N_VGND_c_698_n 0.00562151f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_46 VNB N_VGND_c_699_n 0.095433f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.492
cc_47 VNB N_VGND_c_700_n 0.0175706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_701_n 0.0188229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_702_n 0.32741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_703_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_704_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_D1_c_105_n 0.0174197f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_53 VPB N_D1_c_106_n 0.0157008f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_54 VPB N_D1_c_103_n 0.0159554f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.492
cc_55 VPB N_C1_c_152_n 0.0158345f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_56 VPB N_C1_c_153_n 0.0157476f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_57 VPB N_C1_c_151_n 0.0132422f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_58 VPB N_B1_c_214_n 0.0159376f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_59 VPB N_B1_c_207_n 0.00805528f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.22
cc_60 VPB N_B1_c_216_n 0.0179811f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_61 VPB N_B1_c_210_n 0.00613405f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.492
cc_62 VPB N_B1_c_211_n 0.0079228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_B1_c_212_n 0.0155439f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_64 VPB B1 0.0117591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A2_c_275_n 0.0184237f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_66 VPB N_A2_c_276_n 0.0147903f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_67 VPB A2 0.00786948f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.492
cc_68 VPB N_A2_c_274_n 0.0200394f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_69 VPB N_A1_c_323_n 0.0157756f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_70 VPB N_A1_c_324_n 0.0212384f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_71 VPB A1 0.0110388f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.492
cc_72 VPB N_A1_c_322_n 0.0247753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_364_n 0.011928f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.492
cc_74 VPB N_VPWR_c_365_n 0.0563437f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_75 VPB N_VPWR_c_366_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_76 VPB N_VPWR_c_367_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_368_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_369_n 0.0149451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_370_n 0.00651803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_371_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_372_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_373_n 0.0389676f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_374_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_363_n 0.0906651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_376_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_377_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_378_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_379_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_Y_c_444_n 0.00652689f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_90 VPB N_Y_c_445_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_91 VPB N_Y_c_446_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_Y_c_447_n 0.0117034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_Y_c_448_n 0.00183152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB Y 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_697_368#_c_529_n 0.00557702f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_96 VPB N_A_697_368#_c_530_n 0.00523584f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.492
cc_97 VPB N_A_697_368#_c_531_n 0.00384138f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.492
cc_98 VPB N_A_697_368#_c_532_n 0.0075506f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_99 VPB N_A_697_368#_c_533_n 0.035396f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_100 N_D1_c_101_n N_C1_M1004_g 0.0120716f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_101 N_D1_c_103_n N_C1_M1004_g 0.0206777f $X=0.99 $Y=1.492 $X2=0 $Y2=0
cc_102 N_D1_c_106_n N_C1_c_152_n 0.0269318f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_103 N_D1_c_103_n C1 0.00147401f $X=0.99 $Y=1.492 $X2=0 $Y2=0
cc_104 N_D1_c_103_n N_C1_c_151_n 0.00555101f $X=0.99 $Y=1.492 $X2=0 $Y2=0
cc_105 N_D1_c_105_n N_VPWR_c_365_n 0.0100892f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_106 N_D1_c_102_n N_VPWR_c_365_n 0.00185549f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_107 D1 N_VPWR_c_365_n 0.0149782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_108 N_D1_c_106_n N_VPWR_c_366_n 0.00750878f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_109 N_D1_c_105_n N_VPWR_c_371_n 0.00445602f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_110 N_D1_c_106_n N_VPWR_c_371_n 0.00445602f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_111 N_D1_c_105_n N_VPWR_c_363_n 0.00861209f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_112 N_D1_c_106_n N_VPWR_c_363_n 0.00857432f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_113 N_D1_c_101_n N_Y_c_450_n 0.00519789f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_114 N_D1_c_106_n N_Y_c_444_n 0.0161261f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_115 N_D1_c_103_n N_Y_c_444_n 6.95666e-19 $X=0.99 $Y=1.492 $X2=0 $Y2=0
cc_116 N_D1_c_106_n N_Y_c_448_n 8.20931e-19 $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_117 N_D1_c_105_n Y 0.00182425f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_118 N_D1_c_106_n Y 0.00103342f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_119 N_D1_c_103_n Y 0.033422f $X=0.99 $Y=1.492 $X2=0 $Y2=0
cc_120 D1 Y 0.0153466f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_121 N_D1_c_105_n Y 0.00304071f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_122 N_D1_c_106_n Y 7.21551e-19 $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_123 N_D1_c_100_n N_Y_c_443_n 0.00446631f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_124 N_D1_c_101_n N_Y_c_443_n 0.0046202f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_125 N_D1_c_103_n N_Y_c_443_n 0.00997992f $X=0.99 $Y=1.492 $X2=0 $Y2=0
cc_126 D1 N_Y_c_443_n 0.0125724f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_127 N_D1_c_105_n Y 0.0118573f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_128 N_D1_c_106_n Y 0.0121613f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_129 N_D1_c_100_n N_A_40_74#_c_568_n 0.00904821f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_130 N_D1_c_101_n N_A_40_74#_c_568_n 6.7158e-19 $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_131 N_D1_c_102_n N_A_40_74#_c_568_n 0.00177966f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_132 D1 N_A_40_74#_c_568_n 0.0219843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_133 N_D1_c_100_n N_A_40_74#_c_569_n 0.0100245f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_134 N_D1_c_101_n N_A_40_74#_c_569_n 0.0120041f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_135 N_D1_c_100_n N_A_40_74#_c_570_n 0.00282152f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_136 N_D1_c_100_n N_VGND_c_699_n 0.00278247f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_137 N_D1_c_101_n N_VGND_c_699_n 0.00278271f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_138 N_D1_c_100_n N_VGND_c_702_n 0.00357287f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_139 N_D1_c_101_n N_VGND_c_702_n 0.00353526f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_140 N_C1_c_153_n N_B1_c_214_n 0.0244004f $X=1.945 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_141 C1 N_B1_c_210_n 4.71864e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_C1_c_151_n N_B1_c_210_n 0.0123196f $X=1.92 $Y=1.532 $X2=0 $Y2=0
cc_143 C1 B1 0.0103841f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_C1_c_151_n B1 0.0044044f $X=1.92 $Y=1.532 $X2=0 $Y2=0
cc_145 N_C1_c_152_n N_VPWR_c_366_n 0.00646055f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_146 N_C1_c_152_n N_VPWR_c_367_n 0.00445602f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_147 N_C1_c_153_n N_VPWR_c_367_n 0.00445602f $X=1.945 $Y=1.765 $X2=0 $Y2=0
cc_148 N_C1_c_153_n N_VPWR_c_368_n 0.00486623f $X=1.945 $Y=1.765 $X2=0 $Y2=0
cc_149 N_C1_c_152_n N_VPWR_c_363_n 0.00858104f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_150 N_C1_c_153_n N_VPWR_c_363_n 0.00857673f $X=1.945 $Y=1.765 $X2=0 $Y2=0
cc_151 N_C1_c_152_n N_Y_c_444_n 0.0132143f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_152 C1 N_Y_c_444_n 0.0153556f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_153 N_C1_c_151_n N_Y_c_444_n 8.8068e-19 $X=1.92 $Y=1.532 $X2=0 $Y2=0
cc_154 N_C1_c_152_n N_Y_c_445_n 0.00997113f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_155 N_C1_c_153_n N_Y_c_445_n 0.0109808f $X=1.945 $Y=1.765 $X2=0 $Y2=0
cc_156 N_C1_c_153_n N_Y_c_471_n 0.0138274f $X=1.945 $Y=1.765 $X2=0 $Y2=0
cc_157 C1 N_Y_c_471_n 0.00561225f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_158 N_C1_c_153_n N_Y_c_446_n 6.45594e-19 $X=1.945 $Y=1.765 $X2=0 $Y2=0
cc_159 N_C1_c_152_n N_Y_c_448_n 0.00420532f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_160 N_C1_c_153_n N_Y_c_448_n 0.00409391f $X=1.945 $Y=1.765 $X2=0 $Y2=0
cc_161 C1 N_Y_c_448_n 0.0280913f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_162 N_C1_c_151_n N_Y_c_448_n 0.00308885f $X=1.92 $Y=1.532 $X2=0 $Y2=0
cc_163 C1 Y 0.0111203f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_164 N_C1_c_151_n Y 9.2209e-19 $X=1.92 $Y=1.532 $X2=0 $Y2=0
cc_165 N_C1_M1004_g N_Y_c_443_n 5.93224e-19 $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_166 C1 N_Y_c_443_n 0.00514333f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_167 N_C1_c_152_n Y 6.39139e-19 $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_168 N_C1_M1004_g N_A_40_74#_c_569_n 9.48753e-19 $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_169 N_C1_M1004_g N_A_40_74#_c_571_n 2.64945e-19 $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_170 N_C1_M1004_g N_A_40_74#_c_572_n 0.00100394f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_171 N_C1_M1005_g N_A_40_74#_c_572_n 0.0104532f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_172 C1 N_A_40_74#_c_572_n 0.003612f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_173 N_C1_c_151_n N_A_40_74#_c_572_n 0.00105246f $X=1.92 $Y=1.532 $X2=0 $Y2=0
cc_174 N_C1_M1004_g N_A_40_74#_c_586_n 0.0106874f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_175 N_C1_M1005_g N_A_40_74#_c_586_n 0.00854195f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_176 C1 N_A_40_74#_c_586_n 0.0319834f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_177 N_C1_c_151_n N_A_40_74#_c_586_n 8.8457e-19 $X=1.92 $Y=1.532 $X2=0 $Y2=0
cc_178 N_C1_M1005_g N_A_299_74#_c_608_n 0.0112994f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_179 N_C1_M1004_g N_A_299_74#_c_609_n 0.00608065f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_180 N_C1_M1005_g N_A_299_74#_c_609_n 4.46617e-19 $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_181 N_C1_M1005_g N_A_510_74#_c_634_n 8.65009e-19 $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_182 N_C1_M1005_g N_A_510_74#_c_636_n 0.00183941f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_183 N_C1_M1004_g N_VGND_c_699_n 0.0043213f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_184 N_C1_M1005_g N_VGND_c_699_n 0.00278271f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_185 N_C1_M1004_g N_VGND_c_702_n 0.00447557f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_186 N_C1_M1005_g N_VGND_c_702_n 0.00359085f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B1_M1009_g N_A2_M1001_g 0.0169057f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_188 B1 N_A2_c_275_n 3.21358e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_189 N_B1_c_212_n A2 2.25782e-19 $X=3.335 $Y=1.515 $X2=0 $Y2=0
cc_190 B1 A2 0.0290778f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_191 N_B1_c_212_n N_A2_c_274_n 0.0169057f $X=3.335 $Y=1.515 $X2=0 $Y2=0
cc_192 B1 N_A2_c_274_n 0.00593555f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_193 N_B1_c_214_n N_VPWR_c_368_n 0.00486623f $X=2.395 $Y=1.765 $X2=0 $Y2=0
cc_194 N_B1_c_216_n N_VPWR_c_369_n 0.00714506f $X=2.845 $Y=1.765 $X2=0 $Y2=0
cc_195 N_B1_c_214_n N_VPWR_c_372_n 0.00445602f $X=2.395 $Y=1.765 $X2=0 $Y2=0
cc_196 N_B1_c_216_n N_VPWR_c_372_n 0.00445602f $X=2.845 $Y=1.765 $X2=0 $Y2=0
cc_197 N_B1_c_214_n N_VPWR_c_363_n 0.00857673f $X=2.395 $Y=1.765 $X2=0 $Y2=0
cc_198 N_B1_c_216_n N_VPWR_c_363_n 0.00862391f $X=2.845 $Y=1.765 $X2=0 $Y2=0
cc_199 N_B1_c_214_n N_Y_c_471_n 0.0156348f $X=2.395 $Y=1.765 $X2=0 $Y2=0
cc_200 N_B1_c_214_n N_Y_c_446_n 0.0103431f $X=2.395 $Y=1.765 $X2=0 $Y2=0
cc_201 N_B1_c_216_n N_Y_c_446_n 0.01498f $X=2.845 $Y=1.765 $X2=0 $Y2=0
cc_202 N_B1_c_216_n N_Y_c_447_n 0.0139279f $X=2.845 $Y=1.765 $X2=0 $Y2=0
cc_203 N_B1_c_211_n N_Y_c_447_n 0.00288932f $X=2.985 $Y=1.515 $X2=0 $Y2=0
cc_204 B1 N_Y_c_447_n 0.0714268f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_205 N_B1_c_214_n N_Y_c_448_n 0.00144253f $X=2.395 $Y=1.765 $X2=0 $Y2=0
cc_206 N_B1_c_214_n N_Y_c_490_n 8.98002e-19 $X=2.395 $Y=1.765 $X2=0 $Y2=0
cc_207 N_B1_c_207_n N_Y_c_490_n 0.00132043f $X=2.755 $Y=1.605 $X2=0 $Y2=0
cc_208 N_B1_c_216_n N_Y_c_490_n 4.27055e-19 $X=2.845 $Y=1.765 $X2=0 $Y2=0
cc_209 B1 N_Y_c_490_n 0.0201879f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_210 N_B1_M1007_g N_A_40_74#_c_572_n 0.00129437f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B1_M1007_g N_A_299_74#_c_608_n 0.0132622f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B1_M1009_g N_A_299_74#_c_608_n 0.00500371f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B1_M1009_g N_A_299_74#_c_615_n 0.00491451f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B1_M1007_g N_A_510_74#_c_634_n 0.00750528f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_215 N_B1_M1009_g N_A_510_74#_c_634_n 8.63392e-19 $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B1_M1007_g N_A_510_74#_c_635_n 0.0093986f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_217 N_B1_M1009_g N_A_510_74#_c_635_n 0.0134662f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_218 N_B1_c_212_n N_A_510_74#_c_635_n 0.00381149f $X=3.335 $Y=1.515 $X2=0
+ $Y2=0
cc_219 B1 N_A_510_74#_c_635_n 0.0512198f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_220 N_B1_c_207_n N_A_510_74#_c_636_n 0.00131159f $X=2.755 $Y=1.605 $X2=0
+ $Y2=0
cc_221 N_B1_M1007_g N_A_510_74#_c_636_n 0.00326704f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B1_c_211_n N_A_510_74#_c_636_n 0.00135494f $X=2.985 $Y=1.515 $X2=0
+ $Y2=0
cc_223 B1 N_A_510_74#_c_636_n 0.0289808f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_224 N_B1_M1009_g N_A_510_74#_c_637_n 3.92031e-19 $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_225 B1 N_A_510_74#_c_638_n 3.67275e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_226 B1 N_A_510_74#_c_642_n 0.0153286f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B1_M1009_g N_VGND_c_697_n 5.13093e-19 $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B1_M1007_g N_VGND_c_699_n 0.00278271f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B1_M1009_g N_VGND_c_699_n 0.00430908f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B1_M1007_g N_VGND_c_702_n 0.00359085f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B1_M1009_g N_VGND_c_702_n 0.00817424f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A2_M1015_g N_A1_M1006_g 0.0195237f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A2_c_276_n N_A1_c_323_n 0.0120519f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_234 A2 A1 0.0273144f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_235 A2 N_A1_c_322_n 0.013055f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_236 N_A2_c_274_n N_A1_c_322_n 0.0205436f $X=4.29 $Y=1.557 $X2=0 $Y2=0
cc_237 N_A2_c_275_n N_VPWR_c_369_n 8.40374e-19 $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A2_c_275_n N_VPWR_c_373_n 0.00278271f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A2_c_276_n N_VPWR_c_373_n 0.00278271f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A2_c_275_n N_VPWR_c_363_n 0.00358624f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A2_c_276_n N_VPWR_c_363_n 0.00353907f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A2_c_275_n N_Y_c_447_n 0.0180205f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A2_c_275_n N_Y_c_495_n 0.0139331f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_244 N_A2_c_276_n N_Y_c_495_n 0.0091595f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_245 A2 N_Y_c_495_n 0.0210582f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A2_c_274_n N_Y_c_495_n 0.00137133f $X=4.29 $Y=1.557 $X2=0 $Y2=0
cc_247 N_A2_c_275_n N_A_697_368#_c_530_n 0.0136093f $X=3.855 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A2_c_276_n N_A_697_368#_c_530_n 0.012504f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_249 A2 N_A_697_368#_c_536_n 0.0150276f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_250 A2 N_A_697_368#_c_537_n 0.00285429f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_251 N_A2_M1001_g N_A_299_74#_c_608_n 3.00542e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A2_M1001_g N_A_510_74#_c_637_n 3.92313e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1001_g N_A_510_74#_c_638_n 0.0177463f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A2_M1015_g N_A_510_74#_c_638_n 0.0136953f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_255 A2 N_A_510_74#_c_638_n 0.0344116f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_256 N_A2_c_274_n N_A_510_74#_c_638_n 0.00343847f $X=4.29 $Y=1.557 $X2=0 $Y2=0
cc_257 N_A2_M1015_g N_A_510_74#_c_639_n 4.03583e-19 $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_258 A2 N_A_510_74#_c_640_n 3.30926e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_259 A2 N_A_510_74#_c_643_n 0.0223224f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_260 N_A2_M1001_g N_VGND_c_697_n 0.0105278f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A2_M1015_g N_VGND_c_697_n 0.0091926f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A2_M1001_g N_VGND_c_699_n 0.00383152f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A2_M1015_g N_VGND_c_700_n 0.00444681f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A2_M1001_g N_VGND_c_702_n 0.00757637f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A2_M1015_g N_VGND_c_702_n 0.00877616f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A1_c_323_n N_VPWR_c_370_n 0.0102822f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A1_c_324_n N_VPWR_c_370_n 0.0068696f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A1_c_323_n N_VPWR_c_373_n 0.00413917f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_269 N_A1_c_324_n N_VPWR_c_374_n 0.00445602f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_270 N_A1_c_323_n N_VPWR_c_363_n 0.0081781f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A1_c_324_n N_VPWR_c_363_n 0.00860873f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A1_c_323_n N_A_697_368#_c_530_n 0.00125031f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A1_c_323_n N_A_697_368#_c_537_n 0.0175092f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_A1_c_324_n N_A_697_368#_c_537_n 0.0122806f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_275 A1 N_A_697_368#_c_537_n 0.0280571f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_276 N_A1_c_322_n N_A_697_368#_c_537_n 0.00334184f $X=5.25 $Y=1.515 $X2=0
+ $Y2=0
cc_277 N_A1_c_324_n N_A_697_368#_c_532_n 4.27055e-19 $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_278 A1 N_A_697_368#_c_532_n 0.0255993f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_279 N_A1_c_322_n N_A_697_368#_c_532_n 3.26146e-19 $X=5.25 $Y=1.515 $X2=0
+ $Y2=0
cc_280 N_A1_c_323_n N_A_697_368#_c_533_n 8.85795e-19 $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A1_c_324_n N_A_697_368#_c_533_n 0.0102401f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A1_M1006_g N_A_510_74#_c_639_n 0.00913563f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A1_M1010_g N_A_510_74#_c_639_n 9.66583e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A1_M1006_g N_A_510_74#_c_640_n 0.0151442f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A1_M1010_g N_A_510_74#_c_640_n 0.0140467f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_286 A1 N_A_510_74#_c_640_n 0.0542669f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_287 N_A1_c_322_n N_A_510_74#_c_640_n 0.00728036f $X=5.25 $Y=1.515 $X2=0 $Y2=0
cc_288 N_A1_M1010_g N_A_510_74#_c_641_n 0.00159319f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A1_M1006_g N_A_510_74#_c_643_n 0.00155819f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A1_M1006_g N_VGND_c_697_n 5.12014e-19 $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A1_M1006_g N_VGND_c_698_n 0.00426511f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A1_M1010_g N_VGND_c_698_n 0.013385f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A1_M1006_g N_VGND_c_700_n 0.00434272f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_294 N_A1_M1010_g N_VGND_c_701_n 0.00383152f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A1_M1006_g N_VGND_c_702_n 0.00820816f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A1_M1010_g N_VGND_c_702_n 0.00761342f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_297 N_VPWR_M1019_s N_Y_c_444_n 0.00275645f $X=1.07 $Y=1.84 $X2=0 $Y2=0
cc_298 N_VPWR_c_366_n N_Y_c_444_n 0.0184684f $X=1.27 $Y=2.305 $X2=0 $Y2=0
cc_299 N_VPWR_c_366_n N_Y_c_445_n 0.0563525f $X=1.27 $Y=2.305 $X2=0 $Y2=0
cc_300 N_VPWR_c_367_n N_Y_c_445_n 0.014552f $X=2.085 $Y=3.33 $X2=0 $Y2=0
cc_301 N_VPWR_c_368_n N_Y_c_445_n 0.0449718f $X=2.17 $Y=2.455 $X2=0 $Y2=0
cc_302 N_VPWR_c_363_n N_Y_c_445_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_303 N_VPWR_M1016_d N_Y_c_471_n 0.00956961f $X=2.02 $Y=1.84 $X2=0 $Y2=0
cc_304 N_VPWR_c_368_n N_Y_c_471_n 0.0136682f $X=2.17 $Y=2.455 $X2=0 $Y2=0
cc_305 N_VPWR_c_368_n N_Y_c_446_n 0.0449718f $X=2.17 $Y=2.455 $X2=0 $Y2=0
cc_306 N_VPWR_c_369_n N_Y_c_446_n 0.0462948f $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_307 N_VPWR_c_372_n N_Y_c_446_n 0.014552f $X=2.985 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_363_n N_Y_c_446_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_M1003_s N_Y_c_447_n 0.00591542f $X=2.92 $Y=1.84 $X2=0 $Y2=0
cc_310 N_VPWR_c_369_n N_Y_c_447_n 0.0202359f $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_311 N_VPWR_c_365_n Y 0.0107081f $X=0.32 $Y=1.985 $X2=0 $Y2=0
cc_312 N_VPWR_c_365_n Y 0.0677182f $X=0.32 $Y=1.985 $X2=0 $Y2=0
cc_313 N_VPWR_c_366_n Y 0.0322767f $X=1.27 $Y=2.305 $X2=0 $Y2=0
cc_314 N_VPWR_c_371_n Y 0.014552f $X=1.105 $Y=3.33 $X2=0 $Y2=0
cc_315 N_VPWR_c_363_n Y 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_316 N_VPWR_c_369_n N_A_697_368#_c_529_n 0.0397233f $X=3.07 $Y=2.455 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_370_n N_A_697_368#_c_530_n 0.0125885f $X=4.98 $Y=2.455 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_373_n N_A_697_368#_c_530_n 0.0582805f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_363_n N_A_697_368#_c_530_n 0.0326824f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_369_n N_A_697_368#_c_531_n 0.0119251f $X=3.07 $Y=2.455 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_373_n N_A_697_368#_c_531_n 0.0179217f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_363_n N_A_697_368#_c_531_n 0.00971942f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_370_n N_A_697_368#_c_555_n 0.040027f $X=4.98 $Y=2.455 $X2=0
+ $Y2=0
cc_324 N_VPWR_M1013_d N_A_697_368#_c_537_n 0.00472015f $X=4.83 $Y=1.84 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_370_n N_A_697_368#_c_537_n 0.0202249f $X=4.98 $Y=2.455 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_370_n N_A_697_368#_c_533_n 0.0266809f $X=4.98 $Y=2.455 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_374_n N_A_697_368#_c_533_n 0.0145938f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_363_n N_A_697_368#_c_533_n 0.0120466f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_329 N_Y_c_447_n N_A_697_368#_M1008_s 0.00660323f $X=3.915 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_330 N_Y_c_447_n N_A_697_368#_c_529_n 0.0202359f $X=3.915 $Y=2.035 $X2=0 $Y2=0
cc_331 N_Y_c_495_n N_A_697_368#_c_529_n 0.0298377f $X=4.08 $Y=2.115 $X2=0 $Y2=0
cc_332 N_Y_M1008_d N_A_697_368#_c_530_n 0.00197722f $X=3.93 $Y=1.84 $X2=0 $Y2=0
cc_333 N_Y_c_495_n N_A_697_368#_c_530_n 0.0160777f $X=4.08 $Y=2.115 $X2=0 $Y2=0
cc_334 N_Y_c_495_n N_A_697_368#_c_536_n 0.013092f $X=4.08 $Y=2.115 $X2=0 $Y2=0
cc_335 N_Y_c_495_n N_A_697_368#_c_555_n 0.039994f $X=4.08 $Y=2.115 $X2=0 $Y2=0
cc_336 N_Y_M1012_s N_A_40_74#_c_569_n 0.00176461f $X=0.635 $Y=0.37 $X2=0 $Y2=0
cc_337 N_Y_c_450_n N_A_40_74#_c_569_n 0.0143448f $X=0.775 $Y=0.86 $X2=0 $Y2=0
cc_338 N_Y_c_444_n N_A_40_74#_c_571_n 0.00549175f $X=1.555 $Y=1.885 $X2=0 $Y2=0
cc_339 N_Y_c_443_n N_A_40_74#_c_571_n 0.00503069f $X=0.77 $Y=1.345 $X2=0 $Y2=0
cc_340 N_A_40_74#_c_586_n N_A_299_74#_M1004_s 0.00470069f $X=1.97 $Y=0.862
+ $X2=-0.19 $Y2=-0.245
cc_341 N_A_40_74#_M1005_d N_A_299_74#_c_608_n 0.00274343f $X=1.995 $Y=0.37 $X2=0
+ $Y2=0
cc_342 N_A_40_74#_c_572_n N_A_299_74#_c_608_n 0.0202288f $X=2.135 $Y=0.86 $X2=0
+ $Y2=0
cc_343 N_A_40_74#_c_586_n N_A_299_74#_c_608_n 0.00364964f $X=1.97 $Y=0.862 $X2=0
+ $Y2=0
cc_344 N_A_40_74#_c_569_n N_A_299_74#_c_609_n 0.0112234f $X=1.12 $Y=0.34 $X2=0
+ $Y2=0
cc_345 N_A_40_74#_c_586_n N_A_299_74#_c_609_n 0.0197079f $X=1.97 $Y=0.862 $X2=0
+ $Y2=0
cc_346 N_A_40_74#_c_572_n N_A_510_74#_c_634_n 0.0286351f $X=2.135 $Y=0.86 $X2=0
+ $Y2=0
cc_347 N_A_40_74#_c_572_n N_A_510_74#_c_636_n 0.00854265f $X=2.135 $Y=0.86 $X2=0
+ $Y2=0
cc_348 N_A_40_74#_c_569_n N_VGND_c_699_n 0.050626f $X=1.12 $Y=0.34 $X2=0 $Y2=0
cc_349 N_A_40_74#_c_570_n N_VGND_c_699_n 0.0235688f $X=0.51 $Y=0.34 $X2=0 $Y2=0
cc_350 N_A_40_74#_c_569_n N_VGND_c_702_n 0.028285f $X=1.12 $Y=0.34 $X2=0 $Y2=0
cc_351 N_A_40_74#_c_570_n N_VGND_c_702_n 0.0127152f $X=0.51 $Y=0.34 $X2=0 $Y2=0
cc_352 N_A_40_74#_c_586_n N_VGND_c_702_n 0.00653179f $X=1.97 $Y=0.862 $X2=0
+ $Y2=0
cc_353 N_A_299_74#_c_608_n N_A_510_74#_M1007_d 0.00273752f $X=3.03 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_354 N_A_299_74#_c_608_n N_A_510_74#_c_634_n 0.0203278f $X=3.03 $Y=0.34 $X2=0
+ $Y2=0
cc_355 N_A_299_74#_M1007_s N_A_510_74#_c_635_n 0.00250873f $X=2.985 $Y=0.37
+ $X2=0 $Y2=0
cc_356 N_A_299_74#_c_608_n N_A_510_74#_c_635_n 0.00304353f $X=3.03 $Y=0.34 $X2=0
+ $Y2=0
cc_357 N_A_299_74#_c_615_n N_A_510_74#_c_635_n 0.0207721f $X=3.195 $Y=0.635
+ $X2=0 $Y2=0
cc_358 N_A_299_74#_c_608_n N_A_510_74#_c_637_n 0.00370621f $X=3.03 $Y=0.34 $X2=0
+ $Y2=0
cc_359 N_A_299_74#_c_608_n N_VGND_c_697_n 0.0029789f $X=3.03 $Y=0.34 $X2=0 $Y2=0
cc_360 N_A_299_74#_c_608_n N_VGND_c_699_n 0.101637f $X=3.03 $Y=0.34 $X2=0 $Y2=0
cc_361 N_A_299_74#_c_609_n N_VGND_c_699_n 0.0225845f $X=1.635 $Y=0.34 $X2=0
+ $Y2=0
cc_362 N_A_299_74#_c_608_n N_VGND_c_702_n 0.0575414f $X=3.03 $Y=0.34 $X2=0 $Y2=0
cc_363 N_A_299_74#_c_609_n N_VGND_c_702_n 0.0124836f $X=1.635 $Y=0.34 $X2=0
+ $Y2=0
cc_364 N_A_510_74#_c_638_n N_VGND_M1001_s 0.00197722f $X=4.42 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_365 N_A_510_74#_c_640_n N_VGND_M1006_s 0.00250873f $X=5.35 $Y=1.095 $X2=0
+ $Y2=0
cc_366 N_A_510_74#_c_637_n N_VGND_c_697_n 0.0182488f $X=3.625 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_A_510_74#_c_638_n N_VGND_c_697_n 0.0172656f $X=4.42 $Y=1.095 $X2=0
+ $Y2=0
cc_368 N_A_510_74#_c_639_n N_VGND_c_697_n 0.0168193f $X=4.505 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_A_510_74#_c_639_n N_VGND_c_698_n 0.0184106f $X=4.505 $Y=0.515 $X2=0
+ $Y2=0
cc_370 N_A_510_74#_c_640_n N_VGND_c_698_n 0.0210288f $X=5.35 $Y=1.095 $X2=0
+ $Y2=0
cc_371 N_A_510_74#_c_641_n N_VGND_c_698_n 0.0182902f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
cc_372 N_A_510_74#_c_637_n N_VGND_c_699_n 0.00749631f $X=3.625 $Y=0.515 $X2=0
+ $Y2=0
cc_373 N_A_510_74#_c_639_n N_VGND_c_700_n 0.0109942f $X=4.505 $Y=0.515 $X2=0
+ $Y2=0
cc_374 N_A_510_74#_c_641_n N_VGND_c_701_n 0.011066f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
cc_375 N_A_510_74#_c_637_n N_VGND_c_702_n 0.0062048f $X=3.625 $Y=0.515 $X2=0
+ $Y2=0
cc_376 N_A_510_74#_c_639_n N_VGND_c_702_n 0.00904371f $X=4.505 $Y=0.515 $X2=0
+ $Y2=0
cc_377 N_A_510_74#_c_641_n N_VGND_c_702_n 0.00915947f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
