* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 a_232_98# GATE_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=2.7852e+12p ps=1.673e+07u
M1001 VGND RESET_B a_1153_74# VNB nlowvt w=740000u l=150000u
+  ad=2.30995e+12p pd=1.387e+07u as=1.776e+11p ps=1.96e+06u
M1002 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.257e+11p pd=2.09e+06u as=0p ps=0u
M1003 a_1153_74# a_670_392# a_913_406# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 VPWR D a_27_136# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1005 VPWR RESET_B a_913_406# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.472e+11p ps=2.86e+06u
M1006 Q a_913_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1007 VGND a_232_98# a_373_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.294e+11p ps=2.1e+06u
M1008 a_586_392# a_27_136# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1009 VPWR a_913_406# a_778_504# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=2.898e+11p ps=2.22e+06u
M1010 Q a_913_406# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1011 VGND a_913_406# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_670_392# a_232_98# a_697_74# VNB nlowvt w=640000u l=150000u
+  ad=1.915e+11p pd=1.93e+06u as=1.536e+11p ps=1.76e+06u
M1013 a_913_406# a_670_392# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_913_406# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_697_74# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_232_98# a_373_82# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1017 a_778_504# a_232_98# a_670_392# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=3.371e+11p ps=2.78e+06u
M1018 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1019 VGND a_913_406# a_870_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1020 a_670_392# a_373_82# a_586_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_870_74# a_373_82# a_670_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
