* File: sky130_fd_sc_hs__a21bo_2.spice
* Created: Thu Aug 27 20:24:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a21bo_2.pex.spice"
.subckt sky130_fd_sc_hs__a21bo_2  VNB VPB B1_N A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_B1_N_M1009_g N_A_32_368#_M1009_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.113368 AS=0.14575 PD=0.959302 PS=1.63 NRD=32.964 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1000 N_VGND_M1009_d N_A_187_244#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.152532 AS=0.1036 PD=1.2907 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_187_244#_M1003_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.24605 AS=0.1036 PD=1.405 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1001 N_A_187_244#_M1001_d N_A_32_368#_M1001_g N_VGND_M1003_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.24605 PD=1.02 PS=1.405 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.8 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 A_587_74# N_A1_M1010_g N_A_187_244#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g A_587_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=17.016 M=1 R=4.93333 SA=75002.7 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_B1_N_M1002_g N_A_32_368#_M1002_s VPB PSHORT L=0.15
+ W=0.84 AD=0.1644 AS=0.231 PD=1.27286 PS=2.23 NRD=32.9975 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1007_d N_A_187_244#_M1007_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2192 PD=1.42 PS=1.69714 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1011 N_X_M1007_d N_A_187_244#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001
+ SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_A_504_392#_M1005_d N_A_32_368#_M1005_g N_A_187_244#_M1005_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_504_392#_M1005_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_504_392#_M1008_d N_A2_M1008_g N_VPWR_M1006_d VPB PSHORT L=0.15 W=1
+ AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__a21bo_2.pxi.spice"
*
.ends
*
*
