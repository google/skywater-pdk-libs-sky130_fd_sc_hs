* NGSPICE file created from sky130_fd_sc_hs__o32a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_564_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.2032e+12p pd=1.144e+07u as=1.5408e+12p ps=1.279e+07u
M1001 a_564_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A1 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_83_256# A3 a_961_392# VPB pshort w=1e+06u l=150000u
+  ad=6.2e+11p pd=5.24e+06u as=8.9e+11p ps=7.78e+06u
M1004 a_83_256# B2 a_534_388# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=7.4e+11p ps=5.48e+06u
M1005 VGND A2 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_534_388# B2 a_83_256# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_961_392# A3 a_83_256# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_83_256# B1 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=0p ps=0u
M1009 VPWR B1 a_534_388# VPB pshort w=1e+06u l=150000u
+  ad=1.8398e+12p pd=1.418e+07u as=0p ps=0u
M1010 a_1234_392# A2 a_961_392# VPB pshort w=1e+06u l=150000u
+  ad=7.9e+11p pd=5.58e+06u as=0p ps=0u
M1011 VGND A3 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_564_74# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_83_256# VGND VNB nlowvt w=740000u l=150000u
+  ad=5.069e+11p pd=4.33e+06u as=0p ps=0u
M1014 VPWR a_83_256# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=8.064e+11p ps=5.92e+06u
M1015 X a_83_256# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_83_256# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_1234_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1234_392# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_83_256# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_961_392# A2 a_1234_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_564_74# B2 a_83_256# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_83_256# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_83_256# B2 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_83_256# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_564_74# B1 a_83_256# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_534_388# B1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_83_256# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

