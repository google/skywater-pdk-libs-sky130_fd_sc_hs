* File: sky130_fd_sc_hs__nand4bb_4.pxi.spice
* Created: Tue Sep  1 20:10:37 2020
* 
x_PM_SKY130_FD_SC_HS__NAND4BB_4%A_N N_A_N_M1019_g N_A_N_c_178_n N_A_N_c_182_n
+ N_A_N_M1025_g N_A_N_c_183_n N_A_N_M1026_g N_A_N_c_184_n A_N N_A_N_c_180_n
+ PM_SKY130_FD_SC_HS__NAND4BB_4%A_N
x_PM_SKY130_FD_SC_HS__NAND4BB_4%B_N N_B_N_M1022_g N_B_N_c_227_n N_B_N_c_228_n
+ N_B_N_c_230_n N_B_N_M1029_g N_B_N_c_231_n N_B_N_M1032_g B_N N_B_N_c_229_n
+ PM_SKY130_FD_SC_HS__NAND4BB_4%B_N
x_PM_SKY130_FD_SC_HS__NAND4BB_4%A_27_114# N_A_27_114#_M1019_s
+ N_A_27_114#_M1025_d N_A_27_114#_c_284_n N_A_27_114#_M1000_g
+ N_A_27_114#_c_300_n N_A_27_114#_M1020_g N_A_27_114#_c_285_n
+ N_A_27_114#_M1005_g N_A_27_114#_c_301_n N_A_27_114#_M1021_g
+ N_A_27_114#_c_286_n N_A_27_114#_M1011_g N_A_27_114#_c_302_n
+ N_A_27_114#_M1027_g N_A_27_114#_M1031_g N_A_27_114#_c_288_n
+ N_A_27_114#_c_289_n N_A_27_114#_c_305_n N_A_27_114#_M1030_g
+ N_A_27_114#_c_290_n N_A_27_114#_c_291_n N_A_27_114#_c_292_n
+ N_A_27_114#_c_307_n N_A_27_114#_c_308_n N_A_27_114#_c_293_n
+ N_A_27_114#_c_309_n N_A_27_114#_c_294_n N_A_27_114#_c_295_n
+ N_A_27_114#_c_296_n N_A_27_114#_c_297_n N_A_27_114#_c_298_n
+ N_A_27_114#_c_299_n PM_SKY130_FD_SC_HS__NAND4BB_4%A_27_114#
x_PM_SKY130_FD_SC_HS__NAND4BB_4%A_232_114# N_A_232_114#_M1022_d
+ N_A_232_114#_M1029_d N_A_232_114#_c_443_n N_A_232_114#_M1002_g
+ N_A_232_114#_c_444_n N_A_232_114#_c_445_n N_A_232_114#_c_454_n
+ N_A_232_114#_M1001_g N_A_232_114#_c_446_n N_A_232_114#_M1007_g
+ N_A_232_114#_c_455_n N_A_232_114#_M1004_g N_A_232_114#_c_447_n
+ N_A_232_114#_M1017_g N_A_232_114#_c_456_n N_A_232_114#_M1033_g
+ N_A_232_114#_c_448_n N_A_232_114#_M1028_g N_A_232_114#_c_457_n
+ N_A_232_114#_M1035_g N_A_232_114#_c_449_n N_A_232_114#_c_459_n
+ N_A_232_114#_c_460_n N_A_232_114#_c_461_n N_A_232_114#_c_462_n
+ N_A_232_114#_c_463_n N_A_232_114#_c_464_n N_A_232_114#_c_450_n
+ N_A_232_114#_c_451_n N_A_232_114#_c_452_n N_A_232_114#_c_467_n
+ N_A_232_114#_c_453_n PM_SKY130_FD_SC_HS__NAND4BB_4%A_232_114#
x_PM_SKY130_FD_SC_HS__NAND4BB_4%C N_C_c_626_n N_C_M1006_g N_C_M1023_g
+ N_C_c_627_n N_C_M1009_g N_C_M1024_g N_C_c_628_n N_C_M1012_g N_C_M1036_g
+ N_C_c_629_n N_C_M1014_g N_C_M1037_g N_C_c_638_p C N_C_c_624_n N_C_c_625_n
+ N_C_c_631_n PM_SKY130_FD_SC_HS__NAND4BB_4%C
x_PM_SKY130_FD_SC_HS__NAND4BB_4%D N_D_M1003_g N_D_c_723_n N_D_M1010_g
+ N_D_M1008_g N_D_c_724_n N_D_M1015_g N_D_M1013_g N_D_c_725_n N_D_M1016_g
+ N_D_c_726_n N_D_M1018_g N_D_M1034_g D D D D N_D_c_722_n
+ PM_SKY130_FD_SC_HS__NAND4BB_4%D
x_PM_SKY130_FD_SC_HS__NAND4BB_4%VPWR N_VPWR_M1025_s N_VPWR_M1026_s
+ N_VPWR_M1032_s N_VPWR_M1021_s N_VPWR_M1030_s N_VPWR_M1004_s N_VPWR_M1035_s
+ N_VPWR_M1009_s N_VPWR_M1014_s N_VPWR_M1015_s N_VPWR_M1018_s N_VPWR_c_804_n
+ N_VPWR_c_805_n N_VPWR_c_806_n N_VPWR_c_807_n N_VPWR_c_808_n N_VPWR_c_809_n
+ N_VPWR_c_810_n N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_813_n N_VPWR_c_814_n
+ N_VPWR_c_815_n N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_818_n N_VPWR_c_819_n
+ N_VPWR_c_820_n N_VPWR_c_821_n N_VPWR_c_822_n VPWR N_VPWR_c_823_n
+ N_VPWR_c_824_n N_VPWR_c_825_n N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n
+ N_VPWR_c_829_n N_VPWR_c_830_n N_VPWR_c_831_n N_VPWR_c_832_n N_VPWR_c_833_n
+ N_VPWR_c_834_n N_VPWR_c_835_n N_VPWR_c_803_n
+ PM_SKY130_FD_SC_HS__NAND4BB_4%VPWR
x_PM_SKY130_FD_SC_HS__NAND4BB_4%Y N_Y_M1000_s N_Y_M1011_s N_Y_M1020_d
+ N_Y_M1027_d N_Y_M1001_d N_Y_M1033_d N_Y_M1006_d N_Y_M1012_d N_Y_M1010_d
+ N_Y_M1016_d N_Y_c_994_n N_Y_c_998_n N_Y_c_1168_p N_Y_c_977_n N_Y_c_980_n
+ N_Y_c_1005_n N_Y_c_981_n N_Y_c_1037_n N_Y_c_978_n N_Y_c_983_n N_Y_c_984_n
+ N_Y_c_985_n N_Y_c_1068_n N_Y_c_986_n N_Y_c_1077_n N_Y_c_987_n N_Y_c_1096_n
+ N_Y_c_1100_n N_Y_c_988_n N_Y_c_1006_n N_Y_c_1008_n N_Y_c_979_n N_Y_c_1014_n
+ N_Y_c_1015_n N_Y_c_989_n N_Y_c_990_n N_Y_c_991_n N_Y_c_1108_n Y Y
+ PM_SKY130_FD_SC_HS__NAND4BB_4%Y
x_PM_SKY130_FD_SC_HS__NAND4BB_4%VGND N_VGND_M1019_d N_VGND_M1003_s
+ N_VGND_M1013_s N_VGND_c_1179_n N_VGND_c_1180_n N_VGND_c_1181_n VGND
+ N_VGND_c_1182_n N_VGND_c_1183_n N_VGND_c_1184_n N_VGND_c_1185_n
+ N_VGND_c_1186_n N_VGND_c_1187_n N_VGND_c_1188_n N_VGND_c_1189_n
+ PM_SKY130_FD_SC_HS__NAND4BB_4%VGND
x_PM_SKY130_FD_SC_HS__NAND4BB_4%A_374_74# N_A_374_74#_M1000_d
+ N_A_374_74#_M1005_d N_A_374_74#_M1031_d N_A_374_74#_M1007_s
+ N_A_374_74#_M1028_s N_A_374_74#_c_1278_n N_A_374_74#_c_1273_n
+ N_A_374_74#_c_1274_n N_A_374_74#_c_1275_n N_A_374_74#_c_1285_n
+ N_A_374_74#_c_1293_n N_A_374_74#_c_1287_n N_A_374_74#_c_1276_n
+ N_A_374_74#_c_1277_n PM_SKY130_FD_SC_HS__NAND4BB_4%A_374_74#
x_PM_SKY130_FD_SC_HS__NAND4BB_4%A_828_74# N_A_828_74#_M1002_d
+ N_A_828_74#_M1017_d N_A_828_74#_M1023_d N_A_828_74#_M1036_d
+ N_A_828_74#_c_1336_n N_A_828_74#_c_1337_n N_A_828_74#_c_1346_n
+ N_A_828_74#_c_1338_n N_A_828_74#_c_1352_n N_A_828_74#_c_1339_n
+ N_A_828_74#_c_1340_n PM_SKY130_FD_SC_HS__NAND4BB_4%A_828_74#
x_PM_SKY130_FD_SC_HS__NAND4BB_4%A_1229_74# N_A_1229_74#_M1023_s
+ N_A_1229_74#_M1024_s N_A_1229_74#_M1037_s N_A_1229_74#_M1008_d
+ N_A_1229_74#_M1034_d N_A_1229_74#_c_1387_n N_A_1229_74#_c_1388_n
+ N_A_1229_74#_c_1389_n N_A_1229_74#_c_1455_n N_A_1229_74#_c_1390_n
+ N_A_1229_74#_c_1391_n N_A_1229_74#_c_1392_n N_A_1229_74#_c_1393_n
+ N_A_1229_74#_c_1394_n N_A_1229_74#_c_1395_n N_A_1229_74#_c_1396_n
+ N_A_1229_74#_c_1397_n N_A_1229_74#_c_1398_n
+ PM_SKY130_FD_SC_HS__NAND4BB_4%A_1229_74#
cc_1 VNB N_A_N_M1019_g 0.0240966f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.94
cc_2 VNB N_A_N_c_178_n 0.0025227f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.895
cc_3 VNB A_N 0.00259701f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_N_c_180_n 0.019833f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_5 VNB N_B_N_M1022_g 0.0287863f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.94
cc_6 VNB N_B_N_c_227_n 0.0109978f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.625
cc_7 VNB N_B_N_c_228_n 0.0112089f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.895
cc_8 VNB N_B_N_c_229_n 0.0255078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_114#_c_284_n 0.0202274f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_10 VNB N_A_27_114#_c_285_n 0.0171674f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.97
cc_11 VNB N_A_27_114#_c_286_n 0.0162336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_114#_M1031_g 0.0203986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_114#_c_288_n 0.0134264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_114#_c_289_n 0.0998072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_114#_c_290_n 0.0152646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_114#_c_291_n 0.0106894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_114#_c_292_n 0.017588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_114#_c_293_n 0.0083148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_114#_c_294_n 0.00921485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_114#_c_295_n 0.00329688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_114#_c_296_n 0.00789124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_114#_c_297_n 0.00448773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_114#_c_298_n 0.00666148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_114#_c_299_n 0.0151739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_232_114#_c_443_n 0.014463f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_26 VNB N_A_232_114#_c_444_n 0.0101878f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.045
cc_27 VNB N_A_232_114#_c_445_n 0.00855598f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.54
cc_28 VNB N_A_232_114#_c_446_n 0.01378f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.97
cc_29 VNB N_A_232_114#_c_447_n 0.014886f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_30 VNB N_A_232_114#_c_448_n 0.018169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_232_114#_c_449_n 0.00531134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_232_114#_c_450_n 0.00398754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_232_114#_c_451_n 6.33398e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_232_114#_c_452_n 0.00179663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_232_114#_c_453_n 0.107262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_C_M1023_g 0.0287149f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.895
cc_37 VNB N_C_M1024_g 0.0209341f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.97
cc_38 VNB N_C_M1036_g 0.0209341f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.615
cc_39 VNB N_C_M1037_g 0.0219074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_C_c_624_n 0.112909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_C_c_625_n 0.00356294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_D_M1003_g 0.0208435f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.94
cc_43 VNB N_D_M1008_g 0.0203469f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.045
cc_44 VNB N_D_M1013_g 0.0212283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_D_M1034_g 0.0305951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB D 0.0148545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_D_c_722_n 0.131365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VPWR_c_803_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_Y_c_977_n 0.00869888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_Y_c_978_n 0.00429846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_Y_c_979_n 0.00334121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_1179_n 0.0215326f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.54
cc_53 VNB N_VGND_c_1180_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.97
cc_54 VNB N_VGND_c_1181_n 0.00568581f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.615
cc_55 VNB N_VGND_c_1182_n 0.0194575f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_56 VNB N_VGND_c_1183_n 0.172757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1184_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1185_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1186_n 0.536444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1187_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1188_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1189_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_374_74#_c_1273_n 0.00323114f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=1.615
cc_64 VNB N_A_374_74#_c_1274_n 0.00611261f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.615
cc_65 VNB N_A_374_74#_c_1275_n 0.00450137f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.615
cc_66 VNB N_A_374_74#_c_1276_n 0.00209585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_374_74#_c_1277_n 0.00332116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_828_74#_c_1336_n 0.00577659f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.97
cc_69 VNB N_A_828_74#_c_1337_n 0.017247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_828_74#_c_1338_n 0.00402487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_828_74#_c_1339_n 0.00129507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_828_74#_c_1340_n 0.00203124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1229_74#_c_1387_n 0.0038712f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_74 VNB N_A_1229_74#_c_1388_n 0.00307486f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=1.615
cc_75 VNB N_A_1229_74#_c_1389_n 0.00477062f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.615
cc_76 VNB N_A_1229_74#_c_1390_n 0.00633334f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.615
cc_77 VNB N_A_1229_74#_c_1391_n 0.00178889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1229_74#_c_1392_n 0.0042577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1229_74#_c_1393_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1229_74#_c_1394_n 0.0125563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1229_74#_c_1395_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1229_74#_c_1396_n 0.00124819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1229_74#_c_1397_n 0.00713895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1229_74#_c_1398_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VPB N_A_N_c_178_n 0.0200471f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.895
cc_86 VPB N_A_N_c_182_n 0.0173383f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_87 VPB N_A_N_c_183_n 0.0151019f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.045
cc_88 VPB N_A_N_c_184_n 0.0332709f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.97
cc_89 VPB A_N 0.00149699f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_90 VPB N_B_N_c_230_n 0.0143161f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_91 VPB N_B_N_c_231_n 0.0165051f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.045
cc_92 VPB N_B_N_c_229_n 0.0549529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_114#_c_300_n 0.017155f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.045
cc_94 VPB N_A_27_114#_c_301_n 0.0148285f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.97
cc_95 VPB N_A_27_114#_c_302_n 0.0144394f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_96 VPB N_A_27_114#_c_288_n 0.0112038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_114#_c_289_n 0.0496391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_27_114#_c_305_n 0.014451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_27_114#_c_292_n 0.0137798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_114#_c_307_n 0.00638155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_114#_c_308_n 0.00860392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_114#_c_309_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_232_114#_c_454_n 0.0152062f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.54
cc_104 VPB N_A_232_114#_c_455_n 0.0159895f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_105 VPB N_A_232_114#_c_456_n 0.0154627f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_106 VPB N_A_232_114#_c_457_n 0.0149634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_232_114#_c_449_n 0.00647559f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_232_114#_c_459_n 5.53256e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_232_114#_c_460_n 5.69477e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_232_114#_c_461_n 0.00243101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_232_114#_c_462_n 0.0037734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_232_114#_c_463_n 0.00267158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_232_114#_c_464_n 0.00310488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_232_114#_c_450_n 0.00224682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_232_114#_c_451_n 2.94218e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_232_114#_c_467_n 0.00336046f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_232_114#_c_453_n 0.0479101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_C_c_626_n 0.0156841f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_119 VPB N_C_c_627_n 0.016227f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_120 VPB N_C_c_628_n 0.0162421f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.97
cc_121 VPB N_C_c_629_n 0.0161941f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_122 VPB N_C_c_624_n 0.0266257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_C_c_631_n 0.00441337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_D_c_723_n 0.0162381f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.625
cc_125 VPB N_D_c_724_n 0.0155117f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.54
cc_126 VPB N_D_c_725_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_D_c_726_n 0.0179811f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_128 VPB D 0.0180587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_D_c_722_n 0.0246703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_804_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_805_n 0.0350406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_806_n 0.00272921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_807_n 0.00915851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_808_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_809_n 0.0159425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_810_n 0.0026822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_811_n 0.0173363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_812_n 0.00505145f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_813_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_814_n 0.00970163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_815_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_816_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_817_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_818_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_819_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_820_n 0.0498694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_821_n 0.0217466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_822_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_823_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_824_n 0.0186092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_825_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_826_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_827_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_828_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_829_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_830_n 0.00600349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_831_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_832_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_833_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_834_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_835_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_803_n 0.111473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_Y_c_980_n 0.00249359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_Y_c_981_n 0.00243101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_Y_c_978_n 0.00252558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_Y_c_983_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_Y_c_984_n 0.00904199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_Y_c_985_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_Y_c_986_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_Y_c_987_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_Y_c_988_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_Y_c_989_n 2.15868e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_Y_c_990_n 0.00183525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_Y_c_991_n 0.00199581f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB Y 0.00295756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 N_A_N_M1019_g N_B_N_M1022_g 0.0265012f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_177 A_N N_B_N_M1022_g 0.00164408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A_N_c_180_n N_B_N_M1022_g 0.00554618f $X=0.605 $Y=1.615 $X2=0 $Y2=0
cc_179 N_A_N_c_178_n N_B_N_c_228_n 0.00554618f $X=0.595 $Y=1.895 $X2=0 $Y2=0
cc_180 N_A_N_c_184_n N_B_N_c_228_n 0.00247434f $X=0.955 $Y=1.97 $X2=0 $Y2=0
cc_181 N_A_N_c_183_n N_B_N_c_230_n 0.014787f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_182 N_A_N_c_178_n N_B_N_c_229_n 0.00378665f $X=0.595 $Y=1.895 $X2=0 $Y2=0
cc_183 N_A_N_c_184_n N_B_N_c_229_n 0.00653697f $X=0.955 $Y=1.97 $X2=0 $Y2=0
cc_184 N_A_N_M1019_g N_A_27_114#_c_290_n 0.00343265f $X=0.495 $Y=0.94 $X2=0
+ $Y2=0
cc_185 N_A_N_M1019_g N_A_27_114#_c_291_n 0.0059338f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_186 N_A_N_M1019_g N_A_27_114#_c_292_n 0.0174929f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_187 N_A_N_c_184_n N_A_27_114#_c_292_n 0.00228669f $X=0.955 $Y=1.97 $X2=0
+ $Y2=0
cc_188 A_N N_A_27_114#_c_292_n 0.0250768f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A_N_c_182_n N_A_27_114#_c_307_n 0.00941062f $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_190 N_A_N_c_183_n N_A_27_114#_c_307_n 8.08589e-19 $X=0.955 $Y=2.045 $X2=0
+ $Y2=0
cc_191 N_A_N_c_184_n N_A_27_114#_c_307_n 0.0154627f $X=0.955 $Y=1.97 $X2=0 $Y2=0
cc_192 A_N N_A_27_114#_c_307_n 0.0283597f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A_N_M1019_g N_A_27_114#_c_293_n 0.010552f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_194 A_N N_A_27_114#_c_293_n 0.00957008f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A_N_c_180_n N_A_27_114#_c_293_n 0.0034161f $X=0.605 $Y=1.615 $X2=0
+ $Y2=0
cc_196 N_A_N_c_182_n N_A_27_114#_c_309_n 0.00625061f $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_197 N_A_N_c_183_n N_A_27_114#_c_309_n 0.0064138f $X=0.955 $Y=2.045 $X2=0
+ $Y2=0
cc_198 N_A_N_M1019_g N_A_27_114#_c_298_n 0.00422341f $X=0.495 $Y=0.94 $X2=0
+ $Y2=0
cc_199 N_A_N_M1019_g N_A_232_114#_c_449_n 5.52452e-19 $X=0.495 $Y=0.94 $X2=0
+ $Y2=0
cc_200 N_A_N_c_178_n N_A_232_114#_c_449_n 0.00266626f $X=0.595 $Y=1.895 $X2=0
+ $Y2=0
cc_201 N_A_N_c_184_n N_A_232_114#_c_449_n 0.00228473f $X=0.955 $Y=1.97 $X2=0
+ $Y2=0
cc_202 A_N N_A_232_114#_c_449_n 0.0174378f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A_N_c_183_n N_A_232_114#_c_460_n 0.00173684f $X=0.955 $Y=2.045 $X2=0
+ $Y2=0
cc_204 N_A_N_M1019_g N_A_232_114#_c_452_n 0.0015097f $X=0.495 $Y=0.94 $X2=0
+ $Y2=0
cc_205 N_A_N_c_182_n N_VPWR_c_805_n 0.0120175f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_206 N_A_N_c_183_n N_VPWR_c_805_n 5.35985e-19 $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_207 N_A_N_c_182_n N_VPWR_c_806_n 5.05588e-19 $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_208 N_A_N_c_183_n N_VPWR_c_806_n 0.0104182f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_209 N_A_N_c_182_n N_VPWR_c_823_n 0.00413917f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_210 N_A_N_c_183_n N_VPWR_c_823_n 0.00413917f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_211 N_A_N_c_182_n N_VPWR_c_803_n 0.00817726f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_212 N_A_N_c_183_n N_VPWR_c_803_n 0.00817726f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_213 N_A_N_M1019_g N_VGND_c_1179_n 0.0014541f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_214 N_A_N_M1019_g N_VGND_c_1182_n 0.00343632f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_215 N_A_N_M1019_g N_VGND_c_1186_n 0.00484898f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_216 N_B_N_c_229_n N_A_27_114#_c_300_n 0.0180761f $X=1.63 $Y=1.715 $X2=0 $Y2=0
cc_217 B_N N_A_27_114#_c_289_n 0.0012495f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_218 N_B_N_c_229_n N_A_27_114#_c_289_n 0.0093909f $X=1.63 $Y=1.715 $X2=0 $Y2=0
cc_219 N_B_N_M1022_g N_A_27_114#_c_290_n 4.97186e-19 $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_220 N_B_N_M1022_g N_A_27_114#_c_291_n 0.00202668f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_221 N_B_N_M1022_g N_A_27_114#_c_293_n 0.017488f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_222 N_B_N_c_229_n N_A_27_114#_c_293_n 0.00415042f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_223 N_B_N_M1022_g N_A_27_114#_c_294_n 0.00403796f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_224 N_B_N_M1022_g N_A_27_114#_c_295_n 5.59728e-19 $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_225 B_N N_A_27_114#_c_295_n 0.0144744f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_226 N_B_N_c_229_n N_A_27_114#_c_295_n 0.00446309f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_227 N_B_N_c_229_n N_A_27_114#_c_296_n 3.13473e-19 $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_228 B_N N_A_27_114#_c_299_n 0.00252998f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_229 N_B_N_c_229_n N_A_27_114#_c_299_n 0.00395855f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_230 N_B_N_M1022_g N_A_232_114#_c_449_n 0.00619912f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_231 N_B_N_c_227_n N_A_232_114#_c_449_n 0.0106382f $X=1.315 $Y=1.58 $X2=0
+ $Y2=0
cc_232 N_B_N_c_228_n N_A_232_114#_c_449_n 0.002803f $X=1.16 $Y=1.58 $X2=0 $Y2=0
cc_233 B_N N_A_232_114#_c_449_n 0.024406f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B_N_c_229_n N_A_232_114#_c_449_n 0.00551972f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_235 N_B_N_c_227_n N_A_232_114#_c_459_n 5.12562e-19 $X=1.315 $Y=1.58 $X2=0
+ $Y2=0
cc_236 N_B_N_c_230_n N_A_232_114#_c_459_n 0.0168064f $X=1.405 $Y=2.045 $X2=0
+ $Y2=0
cc_237 B_N N_A_232_114#_c_459_n 0.0246279f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_238 N_B_N_c_229_n N_A_232_114#_c_459_n 0.008331f $X=1.63 $Y=1.715 $X2=0 $Y2=0
cc_239 N_B_N_c_230_n N_A_232_114#_c_461_n 9.00673e-19 $X=1.405 $Y=2.045 $X2=0
+ $Y2=0
cc_240 N_B_N_c_231_n N_A_232_114#_c_461_n 0.0156215f $X=1.855 $Y=2.045 $X2=0
+ $Y2=0
cc_241 N_B_N_c_229_n N_A_232_114#_c_462_n 0.00292018f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_242 B_N N_A_232_114#_c_464_n 0.0134925f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_243 N_B_N_c_229_n N_A_232_114#_c_464_n 0.00234052f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_244 N_B_N_M1022_g N_A_232_114#_c_452_n 0.00790561f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_245 N_B_N_c_227_n N_A_232_114#_c_452_n 0.00601966f $X=1.315 $Y=1.58 $X2=0
+ $Y2=0
cc_246 N_B_N_c_231_n N_A_232_114#_c_467_n 0.0147435f $X=1.855 $Y=2.045 $X2=0
+ $Y2=0
cc_247 N_B_N_c_229_n N_A_232_114#_c_467_n 4.52854e-19 $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_248 N_B_N_c_230_n N_VPWR_c_806_n 0.00970826f $X=1.405 $Y=2.045 $X2=0 $Y2=0
cc_249 N_B_N_c_231_n N_VPWR_c_806_n 5.72226e-19 $X=1.855 $Y=2.045 $X2=0 $Y2=0
cc_250 N_B_N_c_231_n N_VPWR_c_807_n 0.00839337f $X=1.855 $Y=2.045 $X2=0 $Y2=0
cc_251 N_B_N_c_230_n N_VPWR_c_824_n 0.00413917f $X=1.405 $Y=2.045 $X2=0 $Y2=0
cc_252 N_B_N_c_231_n N_VPWR_c_824_n 0.00445602f $X=1.855 $Y=2.045 $X2=0 $Y2=0
cc_253 N_B_N_c_230_n N_VPWR_c_803_n 0.00817726f $X=1.405 $Y=2.045 $X2=0 $Y2=0
cc_254 N_B_N_c_231_n N_VPWR_c_803_n 0.00859819f $X=1.855 $Y=2.045 $X2=0 $Y2=0
cc_255 N_B_N_c_231_n Y 8.96035e-19 $X=1.855 $Y=2.045 $X2=0 $Y2=0
cc_256 N_B_N_M1022_g N_VGND_c_1179_n 0.0014541f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_257 N_B_N_M1022_g N_VGND_c_1183_n 0.00344918f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_258 N_B_N_M1022_g N_VGND_c_1186_n 0.00484898f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_259 N_A_27_114#_c_293_n N_A_232_114#_M1022_d 0.00909254f $X=1.59 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_260 N_A_27_114#_M1031_g N_A_232_114#_c_443_n 0.0160597f $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_261 N_A_27_114#_c_288_n N_A_232_114#_c_445_n 0.00449572f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_262 N_A_27_114#_c_289_n N_A_232_114#_c_445_n 0.0160597f $X=3.71 $Y=1.65 $X2=0
+ $Y2=0
cc_263 N_A_27_114#_c_305_n N_A_232_114#_c_454_n 0.0268074f $X=3.975 $Y=1.765
+ $X2=0 $Y2=0
cc_264 N_A_27_114#_c_307_n N_A_232_114#_c_449_n 0.00509936f $X=0.645 $Y=2.035
+ $X2=0 $Y2=0
cc_265 N_A_27_114#_c_295_n N_A_232_114#_c_449_n 0.00287569f $X=1.76 $Y=1.295
+ $X2=0 $Y2=0
cc_266 N_A_27_114#_c_307_n N_A_232_114#_c_460_n 0.00431295f $X=0.645 $Y=2.035
+ $X2=0 $Y2=0
cc_267 N_A_27_114#_c_309_n N_A_232_114#_c_460_n 0.00519353f $X=0.73 $Y=2.265
+ $X2=0 $Y2=0
cc_268 N_A_27_114#_c_300_n N_A_232_114#_c_462_n 0.00293779f $X=2.575 $Y=1.765
+ $X2=0 $Y2=0
cc_269 N_A_27_114#_c_300_n N_A_232_114#_c_463_n 0.00862797f $X=2.575 $Y=1.765
+ $X2=0 $Y2=0
cc_270 N_A_27_114#_c_301_n N_A_232_114#_c_463_n 0.00710454f $X=3.075 $Y=1.765
+ $X2=0 $Y2=0
cc_271 N_A_27_114#_c_302_n N_A_232_114#_c_463_n 0.00686709f $X=3.525 $Y=1.765
+ $X2=0 $Y2=0
cc_272 N_A_27_114#_c_288_n N_A_232_114#_c_463_n 0.0106376f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_273 N_A_27_114#_c_289_n N_A_232_114#_c_463_n 0.0551803f $X=3.71 $Y=1.65 $X2=0
+ $Y2=0
cc_274 N_A_27_114#_c_305_n N_A_232_114#_c_463_n 0.00613655f $X=3.975 $Y=1.765
+ $X2=0 $Y2=0
cc_275 N_A_27_114#_c_296_n N_A_232_114#_c_463_n 0.0722626f $X=2.495 $Y=1.38
+ $X2=0 $Y2=0
cc_276 N_A_27_114#_c_299_n N_A_232_114#_c_463_n 8.85762e-19 $X=2.155 $Y=1.38
+ $X2=0 $Y2=0
cc_277 N_A_27_114#_c_299_n N_A_232_114#_c_464_n 0.0083714f $X=2.155 $Y=1.38
+ $X2=0 $Y2=0
cc_278 N_A_27_114#_c_288_n N_A_232_114#_c_450_n 0.00366867f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_279 N_A_27_114#_c_289_n N_A_232_114#_c_450_n 0.00275733f $X=3.71 $Y=1.65
+ $X2=0 $Y2=0
cc_280 N_A_27_114#_c_293_n N_A_232_114#_c_452_n 0.0179756f $X=1.59 $Y=0.745
+ $X2=0 $Y2=0
cc_281 N_A_27_114#_c_294_n N_A_232_114#_c_452_n 0.0161513f $X=1.675 $Y=1.21
+ $X2=0 $Y2=0
cc_282 N_A_27_114#_c_295_n N_A_232_114#_c_452_n 0.0103428f $X=1.76 $Y=1.295
+ $X2=0 $Y2=0
cc_283 N_A_27_114#_c_300_n N_A_232_114#_c_467_n 0.00161301f $X=2.575 $Y=1.765
+ $X2=0 $Y2=0
cc_284 N_A_27_114#_c_299_n N_A_232_114#_c_467_n 0.00446079f $X=2.155 $Y=1.38
+ $X2=0 $Y2=0
cc_285 N_A_27_114#_c_288_n N_A_232_114#_c_453_n 0.00857869f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_286 N_A_27_114#_c_289_n N_A_232_114#_c_453_n 0.00500626f $X=3.71 $Y=1.65
+ $X2=0 $Y2=0
cc_287 N_A_27_114#_c_308_n N_VPWR_M1025_s 0.00149394f $X=0.27 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_27_114#_c_307_n N_VPWR_c_805_n 0.0116586f $X=0.645 $Y=2.035 $X2=0
+ $Y2=0
cc_289 N_A_27_114#_c_308_n N_VPWR_c_805_n 0.0139521f $X=0.27 $Y=2.035 $X2=0
+ $Y2=0
cc_290 N_A_27_114#_c_309_n N_VPWR_c_805_n 0.0449718f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_291 N_A_27_114#_c_309_n N_VPWR_c_806_n 0.0384581f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_292 N_A_27_114#_c_300_n N_VPWR_c_807_n 0.00802643f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A_27_114#_c_289_n N_VPWR_c_807_n 9.12666e-19 $X=3.71 $Y=1.65 $X2=0
+ $Y2=0
cc_294 N_A_27_114#_c_300_n N_VPWR_c_808_n 6.24912e-19 $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_27_114#_c_301_n N_VPWR_c_808_n 0.00961101f $X=3.075 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A_27_114#_c_302_n N_VPWR_c_808_n 0.00942577f $X=3.525 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A_27_114#_c_305_n N_VPWR_c_808_n 4.50826e-19 $X=3.975 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A_27_114#_c_302_n N_VPWR_c_809_n 0.00413917f $X=3.525 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_27_114#_c_305_n N_VPWR_c_809_n 0.00413917f $X=3.975 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A_27_114#_c_302_n N_VPWR_c_810_n 4.50826e-19 $X=3.525 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_27_114#_c_305_n N_VPWR_c_810_n 0.00938655f $X=3.975 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_27_114#_c_300_n N_VPWR_c_821_n 0.00319845f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A_27_114#_c_301_n N_VPWR_c_821_n 0.00413917f $X=3.075 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_27_114#_c_309_n N_VPWR_c_823_n 0.00749631f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_305 N_A_27_114#_c_300_n N_VPWR_c_803_n 0.00456434f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_27_114#_c_301_n N_VPWR_c_803_n 0.00818187f $X=3.075 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_27_114#_c_302_n N_VPWR_c_803_n 0.00817726f $X=3.525 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_A_27_114#_c_305_n N_VPWR_c_803_n 0.00817726f $X=3.975 $Y=1.765 $X2=0
+ $Y2=0
cc_309 N_A_27_114#_c_309_n N_VPWR_c_803_n 0.0062048f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_310 N_A_27_114#_c_285_n N_Y_c_994_n 0.0108071f $X=2.765 $Y=1.22 $X2=0 $Y2=0
cc_311 N_A_27_114#_c_286_n N_Y_c_994_n 0.0131525f $X=3.205 $Y=1.22 $X2=0 $Y2=0
cc_312 N_A_27_114#_c_289_n N_Y_c_994_n 7.47057e-19 $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_313 N_A_27_114#_c_297_n N_Y_c_994_n 0.0334364f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_314 N_A_27_114#_c_301_n N_Y_c_998_n 0.0151589f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A_27_114#_c_302_n N_Y_c_998_n 0.0126853f $X=3.525 $Y=1.765 $X2=0 $Y2=0
cc_316 N_A_27_114#_c_289_n N_Y_c_998_n 0.0011308f $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_317 N_A_27_114#_M1031_g N_Y_c_977_n 0.0126146f $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_27_114#_c_288_n N_Y_c_977_n 0.00602266f $X=3.885 $Y=1.65 $X2=0 $Y2=0
cc_319 N_A_27_114#_c_302_n N_Y_c_980_n 2.29968e-19 $X=3.525 $Y=1.765 $X2=0 $Y2=0
cc_320 N_A_27_114#_c_305_n N_Y_c_980_n 2.29968e-19 $X=3.975 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A_27_114#_c_305_n N_Y_c_1005_n 0.0126342f $X=3.975 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A_27_114#_c_289_n N_Y_c_1006_n 0.00152005f $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_323 N_A_27_114#_c_296_n N_Y_c_1006_n 0.0251547f $X=2.495 $Y=1.38 $X2=0 $Y2=0
cc_324 N_A_27_114#_c_300_n N_Y_c_1008_n 0.00568675f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_325 N_A_27_114#_c_289_n N_Y_c_1008_n 0.00144974f $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_326 N_A_27_114#_c_286_n N_Y_c_979_n 0.00303208f $X=3.205 $Y=1.22 $X2=0 $Y2=0
cc_327 N_A_27_114#_M1031_g N_Y_c_979_n 3.32495e-19 $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A_27_114#_c_289_n N_Y_c_979_n 0.00333431f $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_329 N_A_27_114#_c_297_n N_Y_c_979_n 0.00387326f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_330 N_A_27_114#_c_289_n N_Y_c_1014_n 0.00113791f $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_331 N_A_27_114#_c_305_n N_Y_c_1015_n 8.89574e-19 $X=3.975 $Y=1.765 $X2=0
+ $Y2=0
cc_332 N_A_27_114#_c_300_n Y 0.0168628f $X=2.575 $Y=1.765 $X2=0 $Y2=0
cc_333 N_A_27_114#_c_301_n Y 0.0041488f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_334 N_A_27_114#_c_293_n N_VGND_M1019_d 0.0124172f $X=1.59 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_335 N_A_27_114#_c_293_n N_VGND_c_1179_n 0.0251972f $X=1.59 $Y=0.745 $X2=0
+ $Y2=0
cc_336 N_A_27_114#_c_290_n N_VGND_c_1182_n 0.00836867f $X=0.272 $Y=0.83 $X2=0
+ $Y2=0
cc_337 N_A_27_114#_c_293_n N_VGND_c_1182_n 0.00241616f $X=1.59 $Y=0.745 $X2=0
+ $Y2=0
cc_338 N_A_27_114#_c_284_n N_VGND_c_1183_n 0.00278271f $X=2.23 $Y=1.22 $X2=0
+ $Y2=0
cc_339 N_A_27_114#_c_285_n N_VGND_c_1183_n 0.00279474f $X=2.765 $Y=1.22 $X2=0
+ $Y2=0
cc_340 N_A_27_114#_c_286_n N_VGND_c_1183_n 0.00279474f $X=3.205 $Y=1.22 $X2=0
+ $Y2=0
cc_341 N_A_27_114#_M1031_g N_VGND_c_1183_n 0.00278247f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_342 N_A_27_114#_c_293_n N_VGND_c_1183_n 0.012862f $X=1.59 $Y=0.745 $X2=0
+ $Y2=0
cc_343 N_A_27_114#_c_284_n N_VGND_c_1186_n 0.00359383f $X=2.23 $Y=1.22 $X2=0
+ $Y2=0
cc_344 N_A_27_114#_c_285_n N_VGND_c_1186_n 0.00353573f $X=2.765 $Y=1.22 $X2=0
+ $Y2=0
cc_345 N_A_27_114#_c_286_n N_VGND_c_1186_n 0.00352618f $X=3.205 $Y=1.22 $X2=0
+ $Y2=0
cc_346 N_A_27_114#_M1031_g N_VGND_c_1186_n 0.00353524f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_347 N_A_27_114#_c_290_n N_VGND_c_1186_n 0.0111107f $X=0.272 $Y=0.83 $X2=0
+ $Y2=0
cc_348 N_A_27_114#_c_293_n N_VGND_c_1186_n 0.0290944f $X=1.59 $Y=0.745 $X2=0
+ $Y2=0
cc_349 N_A_27_114#_c_293_n N_A_374_74#_c_1278_n 0.0141315f $X=1.59 $Y=0.745
+ $X2=0 $Y2=0
cc_350 N_A_27_114#_c_294_n N_A_374_74#_c_1278_n 0.015495f $X=1.675 $Y=1.21 $X2=0
+ $Y2=0
cc_351 N_A_27_114#_c_299_n N_A_374_74#_c_1278_n 0.013847f $X=2.155 $Y=1.38 $X2=0
+ $Y2=0
cc_352 N_A_27_114#_c_284_n N_A_374_74#_c_1273_n 0.0144073f $X=2.23 $Y=1.22 $X2=0
+ $Y2=0
cc_353 N_A_27_114#_c_285_n N_A_374_74#_c_1273_n 0.00879331f $X=2.765 $Y=1.22
+ $X2=0 $Y2=0
cc_354 N_A_27_114#_c_286_n N_A_374_74#_c_1275_n 0.00818292f $X=3.205 $Y=1.22
+ $X2=0 $Y2=0
cc_355 N_A_27_114#_M1031_g N_A_374_74#_c_1275_n 0.0102111f $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_356 N_A_27_114#_c_286_n N_A_374_74#_c_1285_n 5.47927e-19 $X=3.205 $Y=1.22
+ $X2=0 $Y2=0
cc_357 N_A_27_114#_M1031_g N_A_374_74#_c_1285_n 0.00468221f $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_358 N_A_27_114#_M1031_g N_A_374_74#_c_1287_n 0.00318514f $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_359 N_A_27_114#_c_284_n N_A_374_74#_c_1276_n 8.87476e-19 $X=2.23 $Y=1.22
+ $X2=0 $Y2=0
cc_360 N_A_27_114#_c_285_n N_A_374_74#_c_1276_n 0.00692257f $X=2.765 $Y=1.22
+ $X2=0 $Y2=0
cc_361 N_A_27_114#_c_286_n N_A_374_74#_c_1276_n 0.00653071f $X=3.205 $Y=1.22
+ $X2=0 $Y2=0
cc_362 N_A_27_114#_M1031_g N_A_374_74#_c_1276_n 6.08651e-19 $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_363 N_A_232_114#_c_457_n N_C_c_626_n 0.0231172f $X=5.825 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_364 N_A_232_114#_c_453_n N_C_c_624_n 0.0147623f $X=5.515 $Y=1.475 $X2=0 $Y2=0
cc_365 N_A_232_114#_c_453_n N_C_c_625_n 7.93442e-19 $X=5.515 $Y=1.475 $X2=0
+ $Y2=0
cc_366 N_A_232_114#_c_460_n N_VPWR_M1026_s 0.00285362f $X=1.295 $Y=2.135 $X2=0
+ $Y2=0
cc_367 N_A_232_114#_c_463_n N_VPWR_M1032_s 0.00594521f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_368 N_A_232_114#_c_467_n N_VPWR_M1032_s 0.00356246f $X=2.05 $Y=2.135 $X2=0
+ $Y2=0
cc_369 N_A_232_114#_c_463_n N_VPWR_M1021_s 0.00198204f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_370 N_A_232_114#_c_463_n N_VPWR_M1030_s 5.22224e-19 $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_371 N_A_232_114#_c_450_n N_VPWR_M1030_s 0.00178606f $X=4.315 $Y=1.555 $X2=0
+ $Y2=0
cc_372 N_A_232_114#_c_459_n N_VPWR_c_806_n 0.00102433f $X=1.515 $Y=2.135 $X2=0
+ $Y2=0
cc_373 N_A_232_114#_c_460_n N_VPWR_c_806_n 0.0133439f $X=1.295 $Y=2.135 $X2=0
+ $Y2=0
cc_374 N_A_232_114#_c_461_n N_VPWR_c_806_n 0.0229093f $X=1.63 $Y=2.265 $X2=0
+ $Y2=0
cc_375 N_A_232_114#_c_461_n N_VPWR_c_807_n 0.0384956f $X=1.63 $Y=2.265 $X2=0
+ $Y2=0
cc_376 N_A_232_114#_c_463_n N_VPWR_c_807_n 0.00739494f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_377 N_A_232_114#_c_467_n N_VPWR_c_807_n 0.0104953f $X=2.05 $Y=2.135 $X2=0
+ $Y2=0
cc_378 N_A_232_114#_c_454_n N_VPWR_c_810_n 0.00955095f $X=4.425 $Y=1.765 $X2=0
+ $Y2=0
cc_379 N_A_232_114#_c_455_n N_VPWR_c_810_n 4.97585e-19 $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_380 N_A_232_114#_c_454_n N_VPWR_c_811_n 0.00413917f $X=4.425 $Y=1.765 $X2=0
+ $Y2=0
cc_381 N_A_232_114#_c_455_n N_VPWR_c_811_n 0.00445602f $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_382 N_A_232_114#_c_455_n N_VPWR_c_812_n 0.00594924f $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_383 N_A_232_114#_c_456_n N_VPWR_c_812_n 0.0128349f $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A_232_114#_c_457_n N_VPWR_c_812_n 5.66383e-19 $X=5.825 $Y=1.765 $X2=0
+ $Y2=0
cc_385 N_A_232_114#_c_456_n N_VPWR_c_813_n 5.77599e-19 $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_386 N_A_232_114#_c_457_n N_VPWR_c_813_n 0.012946f $X=5.825 $Y=1.765 $X2=0
+ $Y2=0
cc_387 N_A_232_114#_c_461_n N_VPWR_c_824_n 0.0123628f $X=1.63 $Y=2.265 $X2=0
+ $Y2=0
cc_388 N_A_232_114#_c_456_n N_VPWR_c_825_n 0.00413917f $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_A_232_114#_c_457_n N_VPWR_c_825_n 0.00413917f $X=5.825 $Y=1.765 $X2=0
+ $Y2=0
cc_390 N_A_232_114#_c_454_n N_VPWR_c_803_n 0.00817726f $X=4.425 $Y=1.765 $X2=0
+ $Y2=0
cc_391 N_A_232_114#_c_455_n N_VPWR_c_803_n 0.00857378f $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_392 N_A_232_114#_c_456_n N_VPWR_c_803_n 0.00817726f $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_393 N_A_232_114#_c_457_n N_VPWR_c_803_n 0.00817726f $X=5.825 $Y=1.765 $X2=0
+ $Y2=0
cc_394 N_A_232_114#_c_461_n N_VPWR_c_803_n 0.0101999f $X=1.63 $Y=2.265 $X2=0
+ $Y2=0
cc_395 N_A_232_114#_c_463_n N_Y_M1020_d 0.00250873f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_396 N_A_232_114#_c_463_n N_Y_M1027_d 0.00197722f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_397 N_A_232_114#_c_463_n N_Y_c_998_n 0.03381f $X=4.145 $Y=1.805 $X2=0 $Y2=0
cc_398 N_A_232_114#_c_443_n N_Y_c_977_n 0.00556262f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_399 N_A_232_114#_c_444_n N_Y_c_977_n 0.00428399f $X=4.335 $Y=1.26 $X2=0 $Y2=0
cc_400 N_A_232_114#_c_445_n N_Y_c_977_n 0.00395324f $X=4.14 $Y=1.26 $X2=0 $Y2=0
cc_401 N_A_232_114#_c_446_n N_Y_c_977_n 0.0055884f $X=4.495 $Y=1.185 $X2=0 $Y2=0
cc_402 N_A_232_114#_c_447_n N_Y_c_977_n 0.00599165f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_403 N_A_232_114#_c_448_n N_Y_c_977_n 0.00646677f $X=5.515 $Y=1.185 $X2=0
+ $Y2=0
cc_404 N_A_232_114#_c_463_n N_Y_c_977_n 0.0208641f $X=4.145 $Y=1.805 $X2=0 $Y2=0
cc_405 N_A_232_114#_c_450_n N_Y_c_977_n 0.0131063f $X=4.315 $Y=1.555 $X2=0 $Y2=0
cc_406 N_A_232_114#_c_451_n N_Y_c_977_n 0.07199f $X=5.18 $Y=1.515 $X2=0 $Y2=0
cc_407 N_A_232_114#_c_453_n N_Y_c_977_n 0.0338638f $X=5.515 $Y=1.475 $X2=0 $Y2=0
cc_408 N_A_232_114#_c_454_n N_Y_c_1005_n 0.0136024f $X=4.425 $Y=1.765 $X2=0
+ $Y2=0
cc_409 N_A_232_114#_c_463_n N_Y_c_1005_n 0.0128932f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_410 N_A_232_114#_c_450_n N_Y_c_1005_n 0.0115881f $X=4.315 $Y=1.555 $X2=0
+ $Y2=0
cc_411 N_A_232_114#_c_451_n N_Y_c_1005_n 0.00567887f $X=5.18 $Y=1.515 $X2=0
+ $Y2=0
cc_412 N_A_232_114#_c_454_n N_Y_c_981_n 2.01613e-19 $X=4.425 $Y=1.765 $X2=0
+ $Y2=0
cc_413 N_A_232_114#_c_455_n N_Y_c_981_n 0.00757732f $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_414 N_A_232_114#_c_455_n N_Y_c_1037_n 0.0133259f $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_A_232_114#_c_456_n N_Y_c_1037_n 0.0142854f $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_416 N_A_232_114#_c_451_n N_Y_c_1037_n 0.0337291f $X=5.18 $Y=1.515 $X2=0 $Y2=0
cc_417 N_A_232_114#_c_453_n N_Y_c_1037_n 0.00911851f $X=5.515 $Y=1.475 $X2=0
+ $Y2=0
cc_418 N_A_232_114#_c_456_n N_Y_c_978_n 0.00128638f $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_419 N_A_232_114#_c_457_n N_Y_c_978_n 0.00128638f $X=5.825 $Y=1.765 $X2=0
+ $Y2=0
cc_420 N_A_232_114#_c_451_n N_Y_c_978_n 0.0188915f $X=5.18 $Y=1.515 $X2=0 $Y2=0
cc_421 N_A_232_114#_c_453_n N_Y_c_978_n 0.0313302f $X=5.515 $Y=1.475 $X2=0 $Y2=0
cc_422 N_A_232_114#_c_456_n N_Y_c_983_n 0.00608423f $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_232_114#_c_457_n N_Y_c_983_n 0.0040695f $X=5.825 $Y=1.765 $X2=0 $Y2=0
cc_424 N_A_232_114#_c_457_n N_Y_c_984_n 0.0167636f $X=5.825 $Y=1.765 $X2=0 $Y2=0
cc_425 N_A_232_114#_c_453_n N_Y_c_984_n 0.00297679f $X=5.515 $Y=1.475 $X2=0
+ $Y2=0
cc_426 N_A_232_114#_c_457_n N_Y_c_985_n 3.0288e-19 $X=5.825 $Y=1.765 $X2=0 $Y2=0
cc_427 N_A_232_114#_c_463_n N_Y_c_1008_n 0.0286803f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_428 N_A_232_114#_c_467_n N_Y_c_1008_n 0.00741583f $X=2.05 $Y=2.135 $X2=0
+ $Y2=0
cc_429 N_A_232_114#_c_463_n N_Y_c_979_n 0.00644065f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_430 N_A_232_114#_c_463_n N_Y_c_1014_n 0.0151326f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_431 N_A_232_114#_c_454_n N_Y_c_1015_n 0.00507563f $X=4.425 $Y=1.765 $X2=0
+ $Y2=0
cc_432 N_A_232_114#_c_455_n N_Y_c_1015_n 0.00459155f $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_433 N_A_232_114#_c_456_n N_Y_c_1015_n 0.00102431f $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_434 N_A_232_114#_c_451_n N_Y_c_1015_n 0.0212472f $X=5.18 $Y=1.515 $X2=0 $Y2=0
cc_435 N_A_232_114#_c_453_n N_Y_c_1015_n 0.0069006f $X=5.515 $Y=1.475 $X2=0
+ $Y2=0
cc_436 N_A_232_114#_c_456_n N_Y_c_989_n 9.01568e-19 $X=5.375 $Y=1.765 $X2=0
+ $Y2=0
cc_437 N_A_232_114#_c_457_n N_Y_c_990_n 5.30685e-19 $X=5.825 $Y=1.765 $X2=0
+ $Y2=0
cc_438 N_A_232_114#_c_443_n N_VGND_c_1183_n 0.00328098f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_439 N_A_232_114#_c_446_n N_VGND_c_1183_n 0.00278271f $X=4.495 $Y=1.185 $X2=0
+ $Y2=0
cc_440 N_A_232_114#_c_447_n N_VGND_c_1183_n 0.00278271f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_441 N_A_232_114#_c_448_n N_VGND_c_1183_n 0.00278271f $X=5.515 $Y=1.185 $X2=0
+ $Y2=0
cc_442 N_A_232_114#_c_443_n N_VGND_c_1186_n 0.00427409f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_443 N_A_232_114#_c_446_n N_VGND_c_1186_n 0.00353428f $X=4.495 $Y=1.185 $X2=0
+ $Y2=0
cc_444 N_A_232_114#_c_447_n N_VGND_c_1186_n 0.00354813f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_445 N_A_232_114#_c_448_n N_VGND_c_1186_n 0.00358903f $X=5.515 $Y=1.185 $X2=0
+ $Y2=0
cc_446 N_A_232_114#_c_443_n N_A_374_74#_c_1275_n 0.00120172f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_447 N_A_232_114#_c_443_n N_A_374_74#_c_1293_n 0.0108788f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_448 N_A_232_114#_c_444_n N_A_374_74#_c_1293_n 5.58977e-19 $X=4.335 $Y=1.26
+ $X2=0 $Y2=0
cc_449 N_A_232_114#_c_446_n N_A_374_74#_c_1293_n 0.00843174f $X=4.495 $Y=1.185
+ $X2=0 $Y2=0
cc_450 N_A_232_114#_c_447_n N_A_374_74#_c_1293_n 0.00923324f $X=4.925 $Y=1.185
+ $X2=0 $Y2=0
cc_451 N_A_232_114#_c_448_n N_A_374_74#_c_1293_n 0.00943004f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_452 N_A_232_114#_c_453_n N_A_374_74#_c_1293_n 0.00197046f $X=5.515 $Y=1.475
+ $X2=0 $Y2=0
cc_453 N_A_232_114#_c_447_n N_A_374_74#_c_1277_n 7.8181e-19 $X=4.925 $Y=1.185
+ $X2=0 $Y2=0
cc_454 N_A_232_114#_c_448_n N_A_374_74#_c_1277_n 0.00496352f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_455 N_A_232_114#_c_453_n N_A_374_74#_c_1277_n 0.00582954f $X=5.515 $Y=1.475
+ $X2=0 $Y2=0
cc_456 N_A_232_114#_c_443_n N_A_828_74#_c_1336_n 0.00517186f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_457 N_A_232_114#_c_446_n N_A_828_74#_c_1336_n 0.0125961f $X=4.495 $Y=1.185
+ $X2=0 $Y2=0
cc_458 N_A_232_114#_c_447_n N_A_828_74#_c_1336_n 0.0163854f $X=4.925 $Y=1.185
+ $X2=0 $Y2=0
cc_459 N_A_232_114#_c_448_n N_A_828_74#_c_1337_n 0.012738f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_460 N_A_232_114#_c_448_n N_A_1229_74#_c_1387_n 0.00200707f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_461 N_A_232_114#_c_448_n N_A_1229_74#_c_1389_n 0.00344265f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_462 N_C_M1037_g N_D_M1003_g 0.0127894f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_463 N_C_c_629_n N_D_c_723_n 0.0292057f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_464 N_C_M1037_g D 7.06418e-19 $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_465 N_C_c_638_p D 0.00894849f $X=7.445 $Y=1.485 $X2=0 $Y2=0
cc_466 N_C_c_624_n D 0.00128401f $X=7.725 $Y=1.542 $X2=0 $Y2=0
cc_467 N_C_c_638_p N_D_c_722_n 0.0010812f $X=7.445 $Y=1.485 $X2=0 $Y2=0
cc_468 N_C_c_624_n N_D_c_722_n 0.0254329f $X=7.725 $Y=1.542 $X2=0 $Y2=0
cc_469 N_C_c_626_n N_VPWR_c_813_n 0.00614834f $X=6.275 $Y=1.765 $X2=0 $Y2=0
cc_470 N_C_c_627_n N_VPWR_c_814_n 0.00737447f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_471 N_C_c_628_n N_VPWR_c_814_n 0.00737447f $X=7.275 $Y=1.765 $X2=0 $Y2=0
cc_472 N_C_c_628_n N_VPWR_c_815_n 0.00445602f $X=7.275 $Y=1.765 $X2=0 $Y2=0
cc_473 N_C_c_629_n N_VPWR_c_815_n 0.00445602f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_474 N_C_c_629_n N_VPWR_c_816_n 0.00534288f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_475 N_C_c_626_n N_VPWR_c_826_n 0.00445602f $X=6.275 $Y=1.765 $X2=0 $Y2=0
cc_476 N_C_c_627_n N_VPWR_c_826_n 0.00445602f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_477 N_C_c_626_n N_VPWR_c_803_n 0.00857673f $X=6.275 $Y=1.765 $X2=0 $Y2=0
cc_478 N_C_c_627_n N_VPWR_c_803_n 0.00857797f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_479 N_C_c_628_n N_VPWR_c_803_n 0.00857797f $X=7.275 $Y=1.765 $X2=0 $Y2=0
cc_480 N_C_c_629_n N_VPWR_c_803_n 0.00858104f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_481 N_C_c_624_n N_Y_c_978_n 0.00104018f $X=7.725 $Y=1.542 $X2=0 $Y2=0
cc_482 N_C_c_625_n N_Y_c_978_n 0.0111225f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_483 N_C_c_626_n N_Y_c_984_n 0.0128992f $X=6.275 $Y=1.765 $X2=0 $Y2=0
cc_484 N_C_c_624_n N_Y_c_984_n 4.09899e-19 $X=7.725 $Y=1.542 $X2=0 $Y2=0
cc_485 N_C_c_625_n N_Y_c_984_n 0.0107679f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_486 N_C_c_626_n N_Y_c_985_n 0.0100691f $X=6.275 $Y=1.765 $X2=0 $Y2=0
cc_487 N_C_c_627_n N_Y_c_985_n 0.0109514f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_488 N_C_c_627_n N_Y_c_1068_n 0.0141278f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_489 N_C_c_628_n N_Y_c_1068_n 0.01318f $X=7.275 $Y=1.765 $X2=0 $Y2=0
cc_490 N_C_c_638_p N_Y_c_1068_n 0.0106804f $X=7.445 $Y=1.485 $X2=0 $Y2=0
cc_491 N_C_c_624_n N_Y_c_1068_n 0.00335449f $X=7.725 $Y=1.542 $X2=0 $Y2=0
cc_492 N_C_c_625_n N_Y_c_1068_n 0.00716966f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_493 N_C_c_631_n N_Y_c_1068_n 0.0179859f $X=7.075 $Y=1.55 $X2=0 $Y2=0
cc_494 N_C_c_627_n N_Y_c_986_n 6.63528e-19 $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_495 N_C_c_628_n N_Y_c_986_n 0.0109514f $X=7.275 $Y=1.765 $X2=0 $Y2=0
cc_496 N_C_c_629_n N_Y_c_986_n 0.0112197f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_497 N_C_c_629_n N_Y_c_1077_n 0.0163125f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_498 N_C_c_624_n N_Y_c_1077_n 0.00112245f $X=7.725 $Y=1.542 $X2=0 $Y2=0
cc_499 N_C_c_629_n N_Y_c_987_n 6.04643e-19 $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_500 N_C_c_626_n N_Y_c_990_n 0.00359546f $X=6.275 $Y=1.765 $X2=0 $Y2=0
cc_501 N_C_c_627_n N_Y_c_990_n 0.00369999f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_502 N_C_c_628_n N_Y_c_990_n 0.00114926f $X=7.275 $Y=1.765 $X2=0 $Y2=0
cc_503 N_C_c_624_n N_Y_c_990_n 0.0079942f $X=7.725 $Y=1.542 $X2=0 $Y2=0
cc_504 N_C_c_625_n N_Y_c_990_n 0.0275347f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_505 N_C_c_627_n N_Y_c_991_n 4.01067e-19 $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_506 N_C_c_628_n N_Y_c_991_n 0.00323586f $X=7.275 $Y=1.765 $X2=0 $Y2=0
cc_507 N_C_c_629_n N_Y_c_991_n 0.00335283f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_508 N_C_c_638_p N_Y_c_991_n 0.0231238f $X=7.445 $Y=1.485 $X2=0 $Y2=0
cc_509 N_C_c_624_n N_Y_c_991_n 0.00819757f $X=7.725 $Y=1.542 $X2=0 $Y2=0
cc_510 N_C_M1037_g N_VGND_c_1180_n 4.98172e-19 $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_511 N_C_M1023_g N_VGND_c_1183_n 0.00278247f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_512 N_C_M1024_g N_VGND_c_1183_n 0.00278247f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_513 N_C_M1036_g N_VGND_c_1183_n 0.00278247f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_514 N_C_M1037_g N_VGND_c_1183_n 0.00430908f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_515 N_C_M1023_g N_VGND_c_1186_n 0.00358425f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_516 N_C_M1024_g N_VGND_c_1186_n 0.00353427f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_517 N_C_M1036_g N_VGND_c_1186_n 0.00353427f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_518 N_C_M1037_g N_VGND_c_1186_n 0.00816766f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_519 N_C_M1023_g N_A_828_74#_c_1337_n 0.00987533f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_520 N_C_M1023_g N_A_828_74#_c_1346_n 0.0104366f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_521 N_C_M1024_g N_A_828_74#_c_1346_n 0.00593684f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_522 N_C_M1036_g N_A_828_74#_c_1346_n 5.63827e-19 $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_523 N_C_M1024_g N_A_828_74#_c_1338_n 0.00783479f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_524 N_C_M1036_g N_A_828_74#_c_1338_n 0.00990232f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_525 N_C_M1037_g N_A_828_74#_c_1338_n 0.00412426f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_526 N_C_M1024_g N_A_828_74#_c_1352_n 5.63827e-19 $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_527 N_C_M1036_g N_A_828_74#_c_1352_n 0.00593684f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_528 N_C_M1037_g N_A_828_74#_c_1352_n 0.00473467f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_529 N_C_M1023_g N_A_828_74#_c_1340_n 0.00206753f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_530 N_C_M1024_g N_A_828_74#_c_1340_n 0.00206753f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_531 N_C_M1023_g N_A_1229_74#_c_1388_n 0.0119006f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_532 N_C_M1024_g N_A_1229_74#_c_1388_n 0.0111242f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_533 N_C_c_624_n N_A_1229_74#_c_1388_n 0.00386698f $X=7.725 $Y=1.542 $X2=0
+ $Y2=0
cc_534 N_C_c_625_n N_A_1229_74#_c_1388_n 0.0510561f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_535 N_C_c_624_n N_A_1229_74#_c_1389_n 0.00502748f $X=7.725 $Y=1.542 $X2=0
+ $Y2=0
cc_536 N_C_c_625_n N_A_1229_74#_c_1389_n 0.0157582f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_537 N_C_M1036_g N_A_1229_74#_c_1390_n 0.011119f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_538 N_C_M1037_g N_A_1229_74#_c_1390_n 0.0170077f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_539 N_C_c_638_p N_A_1229_74#_c_1390_n 0.0275868f $X=7.445 $Y=1.485 $X2=0
+ $Y2=0
cc_540 N_C_c_624_n N_A_1229_74#_c_1390_n 0.00234038f $X=7.725 $Y=1.542 $X2=0
+ $Y2=0
cc_541 N_C_M1037_g N_A_1229_74#_c_1391_n 3.92031e-19 $X=7.795 $Y=0.74 $X2=0
+ $Y2=0
cc_542 N_C_c_624_n N_A_1229_74#_c_1396_n 0.00233344f $X=7.725 $Y=1.542 $X2=0
+ $Y2=0
cc_543 N_C_c_631_n N_A_1229_74#_c_1396_n 0.0140843f $X=7.075 $Y=1.55 $X2=0 $Y2=0
cc_544 N_D_c_723_n N_VPWR_c_816_n 0.00671059f $X=8.225 $Y=1.765 $X2=0 $Y2=0
cc_545 N_D_c_723_n N_VPWR_c_817_n 0.00445602f $X=8.225 $Y=1.765 $X2=0 $Y2=0
cc_546 N_D_c_724_n N_VPWR_c_817_n 0.00445602f $X=8.675 $Y=1.765 $X2=0 $Y2=0
cc_547 N_D_c_724_n N_VPWR_c_818_n 0.00486623f $X=8.675 $Y=1.765 $X2=0 $Y2=0
cc_548 N_D_c_725_n N_VPWR_c_818_n 0.00486623f $X=9.125 $Y=1.765 $X2=0 $Y2=0
cc_549 N_D_c_726_n N_VPWR_c_820_n 0.00831454f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_550 D N_VPWR_c_820_n 0.0213189f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_551 N_D_c_722_n N_VPWR_c_820_n 0.00118392f $X=9.585 $Y=1.532 $X2=0 $Y2=0
cc_552 N_D_c_725_n N_VPWR_c_827_n 0.00445602f $X=9.125 $Y=1.765 $X2=0 $Y2=0
cc_553 N_D_c_726_n N_VPWR_c_827_n 0.00445602f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_554 N_D_c_723_n N_VPWR_c_803_n 0.00857432f $X=8.225 $Y=1.765 $X2=0 $Y2=0
cc_555 N_D_c_724_n N_VPWR_c_803_n 0.00857589f $X=8.675 $Y=1.765 $X2=0 $Y2=0
cc_556 N_D_c_725_n N_VPWR_c_803_n 0.00857589f $X=9.125 $Y=1.765 $X2=0 $Y2=0
cc_557 N_D_c_726_n N_VPWR_c_803_n 0.00861084f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_558 N_D_c_723_n N_Y_c_986_n 6.99794e-19 $X=8.225 $Y=1.765 $X2=0 $Y2=0
cc_559 N_D_c_723_n N_Y_c_1077_n 0.0157322f $X=8.225 $Y=1.765 $X2=0 $Y2=0
cc_560 D N_Y_c_1077_n 0.00143862f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_561 N_D_c_723_n N_Y_c_987_n 0.0100939f $X=8.225 $Y=1.765 $X2=0 $Y2=0
cc_562 N_D_c_724_n N_Y_c_987_n 0.0103431f $X=8.675 $Y=1.765 $X2=0 $Y2=0
cc_563 N_D_c_725_n N_Y_c_987_n 6.45594e-19 $X=9.125 $Y=1.765 $X2=0 $Y2=0
cc_564 N_D_c_724_n N_Y_c_1096_n 0.0120074f $X=8.675 $Y=1.765 $X2=0 $Y2=0
cc_565 N_D_c_725_n N_Y_c_1096_n 0.0120074f $X=9.125 $Y=1.765 $X2=0 $Y2=0
cc_566 D N_Y_c_1096_n 0.0397842f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_567 N_D_c_722_n N_Y_c_1096_n 0.00117042f $X=9.585 $Y=1.532 $X2=0 $Y2=0
cc_568 N_D_c_725_n N_Y_c_1100_n 4.27055e-19 $X=9.125 $Y=1.765 $X2=0 $Y2=0
cc_569 N_D_c_726_n N_Y_c_1100_n 0.00203651f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_570 D N_Y_c_1100_n 0.0239985f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_571 N_D_c_722_n N_Y_c_1100_n 0.00129563f $X=9.585 $Y=1.532 $X2=0 $Y2=0
cc_572 N_D_c_724_n N_Y_c_988_n 6.45594e-19 $X=8.675 $Y=1.765 $X2=0 $Y2=0
cc_573 N_D_c_725_n N_Y_c_988_n 0.0103431f $X=9.125 $Y=1.765 $X2=0 $Y2=0
cc_574 N_D_c_726_n N_Y_c_988_n 0.00960826f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_575 N_D_c_723_n N_Y_c_991_n 6.04745e-19 $X=8.225 $Y=1.765 $X2=0 $Y2=0
cc_576 N_D_c_723_n N_Y_c_1108_n 4.27055e-19 $X=8.225 $Y=1.765 $X2=0 $Y2=0
cc_577 N_D_c_724_n N_Y_c_1108_n 4.27055e-19 $X=8.675 $Y=1.765 $X2=0 $Y2=0
cc_578 D N_Y_c_1108_n 0.0239985f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_579 N_D_c_722_n N_Y_c_1108_n 0.00129124f $X=9.585 $Y=1.532 $X2=0 $Y2=0
cc_580 N_D_M1003_g N_VGND_c_1180_n 0.0092592f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_581 N_D_M1008_g N_VGND_c_1180_n 0.00921026f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_582 N_D_M1013_g N_VGND_c_1180_n 4.56715e-19 $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_583 N_D_M1008_g N_VGND_c_1181_n 4.56715e-19 $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_584 N_D_M1013_g N_VGND_c_1181_n 0.00921984f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_585 N_D_M1034_g N_VGND_c_1181_n 0.0054497f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_586 N_D_M1003_g N_VGND_c_1183_n 0.00383152f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_587 N_D_M1008_g N_VGND_c_1184_n 0.00383152f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_588 N_D_M1013_g N_VGND_c_1184_n 0.00383152f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_589 N_D_M1034_g N_VGND_c_1185_n 0.00434272f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_590 N_D_M1003_g N_VGND_c_1186_n 0.00757637f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_591 N_D_M1008_g N_VGND_c_1186_n 0.0075754f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_592 N_D_M1013_g N_VGND_c_1186_n 0.0075754f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_593 N_D_M1034_g N_VGND_c_1186_n 0.00824376f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_594 N_D_M1003_g N_A_828_74#_c_1338_n 3.00542e-19 $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_595 N_D_M1003_g N_A_1229_74#_c_1391_n 3.92313e-19 $X=8.225 $Y=0.74 $X2=0
+ $Y2=0
cc_596 N_D_M1003_g N_A_1229_74#_c_1392_n 0.0159972f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_597 N_D_M1008_g N_A_1229_74#_c_1392_n 0.0124847f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_598 D N_A_1229_74#_c_1392_n 0.0395058f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_599 N_D_c_722_n N_A_1229_74#_c_1392_n 0.00269913f $X=9.585 $Y=1.532 $X2=0
+ $Y2=0
cc_600 N_D_M1008_g N_A_1229_74#_c_1393_n 3.92313e-19 $X=8.655 $Y=0.74 $X2=0
+ $Y2=0
cc_601 N_D_M1013_g N_A_1229_74#_c_1393_n 3.92313e-19 $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_602 N_D_M1013_g N_A_1229_74#_c_1394_n 0.0128832f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_603 N_D_M1034_g N_A_1229_74#_c_1394_n 0.0126756f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_604 D N_A_1229_74#_c_1394_n 0.0792081f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_605 N_D_c_722_n N_A_1229_74#_c_1394_n 0.0101096f $X=9.585 $Y=1.532 $X2=0
+ $Y2=0
cc_606 N_D_M1013_g N_A_1229_74#_c_1395_n 9.27941e-19 $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_607 N_D_M1034_g N_A_1229_74#_c_1395_n 0.00959678f $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_608 N_D_M1003_g N_A_1229_74#_c_1397_n 6.32871e-19 $X=8.225 $Y=0.74 $X2=0
+ $Y2=0
cc_609 D N_A_1229_74#_c_1398_n 0.0147161f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_610 N_D_c_722_n N_A_1229_74#_c_1398_n 0.00232957f $X=9.585 $Y=1.532 $X2=0
+ $Y2=0
cc_611 N_VPWR_M1021_s N_Y_c_998_n 0.00363646f $X=3.15 $Y=1.84 $X2=0 $Y2=0
cc_612 N_VPWR_c_808_n N_Y_c_998_n 0.0171814f $X=3.3 $Y=2.495 $X2=0 $Y2=0
cc_613 N_VPWR_c_808_n N_Y_c_980_n 0.0232805f $X=3.3 $Y=2.495 $X2=0 $Y2=0
cc_614 N_VPWR_c_809_n N_Y_c_980_n 0.0105983f $X=4.035 $Y=3.33 $X2=0 $Y2=0
cc_615 N_VPWR_c_810_n N_Y_c_980_n 0.0232805f $X=4.2 $Y=2.495 $X2=0 $Y2=0
cc_616 N_VPWR_c_803_n N_Y_c_980_n 0.00847107f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_617 N_VPWR_M1030_s N_Y_c_1005_n 0.00393416f $X=4.05 $Y=1.84 $X2=0 $Y2=0
cc_618 N_VPWR_c_810_n N_Y_c_1005_n 0.0171f $X=4.2 $Y=2.495 $X2=0 $Y2=0
cc_619 N_VPWR_c_810_n N_Y_c_981_n 0.022534f $X=4.2 $Y=2.495 $X2=0 $Y2=0
cc_620 N_VPWR_c_811_n N_Y_c_981_n 0.0123628f $X=4.985 $Y=3.33 $X2=0 $Y2=0
cc_621 N_VPWR_c_803_n N_Y_c_981_n 0.0101999f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_622 N_VPWR_M1004_s N_Y_c_1037_n 0.00448384f $X=4.95 $Y=1.84 $X2=0 $Y2=0
cc_623 N_VPWR_c_812_n N_Y_c_1037_n 0.0202249f $X=5.15 $Y=2.355 $X2=0 $Y2=0
cc_624 N_VPWR_c_812_n N_Y_c_983_n 0.0514854f $X=5.15 $Y=2.355 $X2=0 $Y2=0
cc_625 N_VPWR_c_813_n N_Y_c_983_n 0.0523143f $X=6.05 $Y=2.325 $X2=0 $Y2=0
cc_626 N_VPWR_c_825_n N_Y_c_983_n 0.00749631f $X=5.885 $Y=3.33 $X2=0 $Y2=0
cc_627 N_VPWR_c_803_n N_Y_c_983_n 0.0062048f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_M1035_s N_Y_c_984_n 0.00222494f $X=5.9 $Y=1.84 $X2=0 $Y2=0
cc_629 N_VPWR_c_813_n N_Y_c_984_n 0.0154248f $X=6.05 $Y=2.325 $X2=0 $Y2=0
cc_630 N_VPWR_c_813_n N_Y_c_985_n 0.0550114f $X=6.05 $Y=2.325 $X2=0 $Y2=0
cc_631 N_VPWR_c_814_n N_Y_c_985_n 0.0266809f $X=7 $Y=2.455 $X2=0 $Y2=0
cc_632 N_VPWR_c_826_n N_Y_c_985_n 0.014552f $X=6.835 $Y=3.33 $X2=0 $Y2=0
cc_633 N_VPWR_c_803_n N_Y_c_985_n 0.0119791f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_634 N_VPWR_M1009_s N_Y_c_1068_n 0.00608585f $X=6.8 $Y=1.84 $X2=0 $Y2=0
cc_635 N_VPWR_c_814_n N_Y_c_1068_n 0.0232685f $X=7 $Y=2.455 $X2=0 $Y2=0
cc_636 N_VPWR_c_814_n N_Y_c_986_n 0.0266809f $X=7 $Y=2.455 $X2=0 $Y2=0
cc_637 N_VPWR_c_815_n N_Y_c_986_n 0.014552f $X=7.865 $Y=3.33 $X2=0 $Y2=0
cc_638 N_VPWR_c_816_n N_Y_c_986_n 0.0462948f $X=7.95 $Y=2.455 $X2=0 $Y2=0
cc_639 N_VPWR_c_803_n N_Y_c_986_n 0.0119791f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_640 N_VPWR_M1014_s N_Y_c_1077_n 0.0114619f $X=7.8 $Y=1.84 $X2=0 $Y2=0
cc_641 N_VPWR_c_816_n N_Y_c_1077_n 0.0184684f $X=7.95 $Y=2.455 $X2=0 $Y2=0
cc_642 N_VPWR_c_816_n N_Y_c_987_n 0.0266484f $X=7.95 $Y=2.455 $X2=0 $Y2=0
cc_643 N_VPWR_c_817_n N_Y_c_987_n 0.014552f $X=8.815 $Y=3.33 $X2=0 $Y2=0
cc_644 N_VPWR_c_818_n N_Y_c_987_n 0.0449718f $X=8.9 $Y=2.455 $X2=0 $Y2=0
cc_645 N_VPWR_c_803_n N_Y_c_987_n 0.0119791f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_646 N_VPWR_M1015_s N_Y_c_1096_n 0.00412199f $X=8.75 $Y=1.84 $X2=0 $Y2=0
cc_647 N_VPWR_c_818_n N_Y_c_1096_n 0.0136682f $X=8.9 $Y=2.455 $X2=0 $Y2=0
cc_648 N_VPWR_c_820_n N_Y_c_1100_n 0.0121024f $X=9.8 $Y=2.115 $X2=0 $Y2=0
cc_649 N_VPWR_c_818_n N_Y_c_988_n 0.0449718f $X=8.9 $Y=2.455 $X2=0 $Y2=0
cc_650 N_VPWR_c_820_n N_Y_c_988_n 0.0576605f $X=9.8 $Y=2.115 $X2=0 $Y2=0
cc_651 N_VPWR_c_827_n N_Y_c_988_n 0.014552f $X=9.715 $Y=3.33 $X2=0 $Y2=0
cc_652 N_VPWR_c_803_n N_Y_c_988_n 0.0119791f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_653 N_VPWR_c_812_n N_Y_c_1015_n 0.0296971f $X=5.15 $Y=2.355 $X2=0 $Y2=0
cc_654 N_VPWR_c_807_n Y 0.0437224f $X=2.17 $Y=2.495 $X2=0 $Y2=0
cc_655 N_VPWR_c_808_n Y 0.0233984f $X=3.3 $Y=2.495 $X2=0 $Y2=0
cc_656 N_VPWR_c_821_n Y 0.0199831f $X=3.135 $Y=3.33 $X2=0 $Y2=0
cc_657 N_VPWR_c_803_n Y 0.015678f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_658 N_Y_c_994_n N_A_374_74#_M1005_d 0.00349797f $X=3.335 $Y=0.955 $X2=0 $Y2=0
cc_659 N_Y_c_977_n N_A_374_74#_M1031_d 0.00176461f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_660 N_Y_c_977_n N_A_374_74#_M1007_s 0.00176891f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_661 N_Y_c_977_n N_A_374_74#_M1028_s 7.73211e-19 $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_662 N_Y_M1000_s N_A_374_74#_c_1273_n 0.00295551f $X=2.305 $Y=0.37 $X2=0 $Y2=0
cc_663 N_Y_c_994_n N_A_374_74#_c_1273_n 0.00404257f $X=3.335 $Y=0.955 $X2=0
+ $Y2=0
cc_664 N_Y_c_1006_n N_A_374_74#_c_1273_n 0.0199719f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_665 N_Y_M1011_s N_A_374_74#_c_1275_n 0.00176461f $X=3.28 $Y=0.37 $X2=0 $Y2=0
cc_666 N_Y_c_994_n N_A_374_74#_c_1275_n 0.00402702f $X=3.335 $Y=0.955 $X2=0
+ $Y2=0
cc_667 N_Y_c_1168_p N_A_374_74#_c_1275_n 0.012613f $X=3.42 $Y=0.87 $X2=0 $Y2=0
cc_668 N_Y_c_977_n N_A_374_74#_c_1275_n 0.00270072f $X=5.515 $Y=1.175 $X2=0
+ $Y2=0
cc_669 N_Y_c_977_n N_A_374_74#_c_1293_n 0.0870842f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_670 N_Y_c_977_n N_A_374_74#_c_1287_n 0.0153817f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_671 N_Y_c_994_n N_A_374_74#_c_1276_n 0.0165533f $X=3.335 $Y=0.955 $X2=0 $Y2=0
cc_672 N_Y_c_977_n N_A_374_74#_c_1277_n 0.00517215f $X=5.515 $Y=1.175 $X2=0
+ $Y2=0
cc_673 N_Y_c_977_n N_A_828_74#_M1002_d 0.00176891f $X=5.515 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_674 N_Y_c_977_n N_A_828_74#_M1017_d 0.00347389f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_675 N_Y_c_977_n N_A_1229_74#_c_1389_n 0.0028602f $X=5.515 $Y=1.175 $X2=0
+ $Y2=0
cc_676 N_Y_c_984_n N_A_1229_74#_c_1389_n 0.0019066f $X=6.335 $Y=1.905 $X2=0
+ $Y2=0
cc_677 N_Y_c_991_n N_A_1229_74#_c_1390_n 0.00169126f $X=7.5 $Y=1.985 $X2=0 $Y2=0
cc_678 N_VGND_c_1183_n N_A_374_74#_c_1273_n 0.045537f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_679 N_VGND_c_1186_n N_A_374_74#_c_1273_n 0.0257922f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_680 N_VGND_c_1183_n N_A_374_74#_c_1274_n 0.0121867f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_681 N_VGND_c_1186_n N_A_374_74#_c_1274_n 0.00660921f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_682 N_VGND_c_1183_n N_A_374_74#_c_1275_n 0.051499f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_683 N_VGND_c_1186_n N_A_374_74#_c_1275_n 0.0285503f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1183_n N_A_374_74#_c_1293_n 0.00197884f $X=8.275 $Y=0 $X2=0
+ $Y2=0
cc_685 N_VGND_c_1186_n N_A_374_74#_c_1293_n 0.00647053f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_686 N_VGND_c_1183_n N_A_374_74#_c_1276_n 0.0226536f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_687 N_VGND_c_1186_n N_A_374_74#_c_1276_n 0.0124411f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_688 N_VGND_c_1183_n N_A_828_74#_c_1336_n 0.159083f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_689 N_VGND_c_1186_n N_A_828_74#_c_1336_n 0.0896859f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_690 N_VGND_c_1180_n N_A_828_74#_c_1338_n 0.0029789f $X=8.44 $Y=0.57 $X2=0
+ $Y2=0
cc_691 N_VGND_c_1183_n N_A_828_74#_c_1338_n 0.0564897f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_692 N_VGND_c_1186_n N_A_828_74#_c_1338_n 0.0313161f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_693 N_VGND_c_1183_n N_A_828_74#_c_1340_n 0.0231282f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_694 N_VGND_c_1186_n N_A_828_74#_c_1340_n 0.0125338f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_695 N_VGND_c_1180_n N_A_1229_74#_c_1391_n 0.0164567f $X=8.44 $Y=0.57 $X2=0
+ $Y2=0
cc_696 N_VGND_c_1183_n N_A_1229_74#_c_1391_n 0.00749631f $X=8.275 $Y=0 $X2=0
+ $Y2=0
cc_697 N_VGND_c_1186_n N_A_1229_74#_c_1391_n 0.0062048f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_698 N_VGND_M1003_s N_A_1229_74#_c_1392_n 0.00176461f $X=8.3 $Y=0.37 $X2=0
+ $Y2=0
cc_699 N_VGND_c_1180_n N_A_1229_74#_c_1392_n 0.0171619f $X=8.44 $Y=0.57 $X2=0
+ $Y2=0
cc_700 N_VGND_c_1180_n N_A_1229_74#_c_1393_n 0.0164567f $X=8.44 $Y=0.57 $X2=0
+ $Y2=0
cc_701 N_VGND_c_1181_n N_A_1229_74#_c_1393_n 0.0164567f $X=9.3 $Y=0.57 $X2=0
+ $Y2=0
cc_702 N_VGND_c_1184_n N_A_1229_74#_c_1393_n 0.00749631f $X=9.135 $Y=0 $X2=0
+ $Y2=0
cc_703 N_VGND_c_1186_n N_A_1229_74#_c_1393_n 0.0062048f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_704 N_VGND_M1013_s N_A_1229_74#_c_1394_n 0.00250873f $X=9.16 $Y=0.37 $X2=0
+ $Y2=0
cc_705 N_VGND_c_1181_n N_A_1229_74#_c_1394_n 0.0210288f $X=9.3 $Y=0.57 $X2=0
+ $Y2=0
cc_706 N_VGND_c_1181_n N_A_1229_74#_c_1395_n 0.0173003f $X=9.3 $Y=0.57 $X2=0
+ $Y2=0
cc_707 N_VGND_c_1185_n N_A_1229_74#_c_1395_n 0.0145639f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_708 N_VGND_c_1186_n N_A_1229_74#_c_1395_n 0.0119984f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_709 N_A_374_74#_c_1293_n N_A_828_74#_M1002_d 0.003292f $X=5.565 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_710 N_A_374_74#_c_1293_n N_A_828_74#_M1017_d 0.0070998f $X=5.565 $Y=0.835
+ $X2=0 $Y2=0
cc_711 N_A_374_74#_M1007_s N_A_828_74#_c_1336_n 0.00171274f $X=4.57 $Y=0.37
+ $X2=0 $Y2=0
cc_712 N_A_374_74#_c_1275_n N_A_828_74#_c_1336_n 0.0119071f $X=3.685 $Y=0.34
+ $X2=0 $Y2=0
cc_713 N_A_374_74#_c_1293_n N_A_828_74#_c_1336_n 0.0708016f $X=5.565 $Y=0.835
+ $X2=0 $Y2=0
cc_714 N_A_374_74#_M1028_s N_A_828_74#_c_1337_n 0.00273752f $X=5.59 $Y=0.37
+ $X2=0 $Y2=0
cc_715 N_A_374_74#_c_1293_n N_A_828_74#_c_1337_n 0.00442249f $X=5.565 $Y=0.835
+ $X2=0 $Y2=0
cc_716 N_A_374_74#_c_1277_n N_A_828_74#_c_1337_n 0.0194173f $X=5.73 $Y=0.715
+ $X2=0 $Y2=0
cc_717 N_A_374_74#_c_1277_n N_A_1229_74#_c_1387_n 0.02146f $X=5.73 $Y=0.715
+ $X2=0 $Y2=0
cc_718 N_A_828_74#_c_1337_n N_A_1229_74#_M1023_s 0.00273752f $X=6.555 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_719 N_A_828_74#_c_1338_n N_A_1229_74#_M1024_s 0.00176461f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
cc_720 N_A_828_74#_c_1337_n N_A_1229_74#_c_1387_n 0.0185632f $X=6.555 $Y=0.34
+ $X2=0 $Y2=0
cc_721 N_A_828_74#_M1023_d N_A_1229_74#_c_1388_n 0.00176461f $X=6.58 $Y=0.37
+ $X2=0 $Y2=0
cc_722 N_A_828_74#_c_1337_n N_A_1229_74#_c_1388_n 0.0031794f $X=6.555 $Y=0.34
+ $X2=0 $Y2=0
cc_723 N_A_828_74#_c_1346_n N_A_1229_74#_c_1388_n 0.0168793f $X=6.72 $Y=0.58
+ $X2=0 $Y2=0
cc_724 N_A_828_74#_c_1338_n N_A_1229_74#_c_1388_n 0.0031794f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
cc_725 N_A_828_74#_c_1338_n N_A_1229_74#_c_1455_n 0.0124395f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
cc_726 N_A_828_74#_M1036_d N_A_1229_74#_c_1390_n 0.00176461f $X=7.44 $Y=0.37
+ $X2=0 $Y2=0
cc_727 N_A_828_74#_c_1338_n N_A_1229_74#_c_1390_n 0.0031794f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
cc_728 N_A_828_74#_c_1352_n N_A_1229_74#_c_1390_n 0.0168793f $X=7.58 $Y=0.58
+ $X2=0 $Y2=0
cc_729 N_A_828_74#_c_1338_n N_A_1229_74#_c_1391_n 0.00370621f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
