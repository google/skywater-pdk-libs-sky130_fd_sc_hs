* File: sky130_fd_sc_hs__einvn_4.pex.spice
* Created: Thu Aug 27 20:44:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__EINVN_4%A_114_74# 1 2 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 28 29 30 31 33 39
c88 39 0 3.83609e-19 $X=1.13 $Y=0.465
c89 22 0 1.82848e-19 $X=2.98 $Y=1.26
c90 8 0 5.82364e-21 $X=1.295 $Y=1.26
r91 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.145 $X2=1.13 $Y2=1.145
r92 41 43 10.4571 $w=7.35e-07 $l=6.3e-07 $layer=LI1_cond $X=0.92 $Y=0.515
+ $X2=0.92 $Y2=1.145
r93 39 44 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=1.13 $Y=0.465
+ $X2=1.13 $Y2=1.145
r94 38 41 0.829932 $w=7.35e-07 $l=5e-08 $layer=LI1_cond $X=0.92 $Y=0.465
+ $X2=0.92 $Y2=0.515
r95 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=0.465 $X2=1.13 $Y2=0.465
r96 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.79 $Y=1.985
+ $X2=0.79 $Y2=2.815
r97 31 43 6.49103 $w=7.35e-07 $l=2.20624e-07 $layer=LI1_cond $X=0.79 $Y=1.31
+ $X2=0.92 $Y2=1.145
r98 31 33 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.79 $Y=1.31
+ $X2=0.79 $Y2=1.985
r99 27 44 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.13 $Y=1.185 $X2=1.13
+ $Y2=1.145
r100 24 26 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.055 $Y=1.185
+ $X2=3.055 $Y2=0.74
r101 23 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.26
+ $X2=2.625 $Y2=1.26
r102 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.98 $Y=1.26
+ $X2=3.055 $Y2=1.185
r103 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.26
+ $X2=2.7 $Y2=1.26
r104 19 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.625 $Y2=1.26
r105 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.625 $Y2=0.74
r106 18 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.26
+ $X2=2.195 $Y2=1.26
r107 17 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.26
+ $X2=2.625 $Y2=1.26
r108 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.26
+ $X2=2.27 $Y2=1.26
r109 14 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.195 $Y2=1.26
r110 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.195 $Y2=0.74
r111 13 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.26
+ $X2=1.765 $Y2=1.26
r112 12 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.26
+ $X2=2.195 $Y2=1.26
r113 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.26
+ $X2=1.84 $Y2=1.26
r114 9 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=1.26
r115 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=0.74
r116 8 27 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.295 $Y=1.26
+ $X2=1.13 $Y2=1.185
r117 7 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.26
+ $X2=1.765 $Y2=1.26
r118 7 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.69 $Y=1.26
+ $X2=1.295 $Y2=1.26
r119 2 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.84 $X2=0.79 $Y2=2.815
r120 2 33 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.84 $X2=0.79 $Y2=1.985
r121 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_4%TE_B 3 5 7 8 10 12 13 15 17 18 20 22 23 25
+ 27 28 29 30 31 35
c95 35 0 5.82364e-21 $X=0.29 $Y=1.465
c96 30 0 1.87728e-19 $X=2.475 $Y=1.67
c97 28 0 1.20768e-19 $X=1.575 $Y=1.67
c98 23 0 1.40151e-19 $X=2.885 $Y=1.65
c99 20 0 9.04372e-20 $X=2.475 $Y=1.765
c100 18 0 1.72388e-19 $X=2.385 $Y=1.65
c101 8 0 1.69662e-19 $X=1.485 $Y=1.65
r102 34 36 17.8697 $w=4.99e-07 $l=1.85e-07 $layer=POLY_cond $X=0.39 $Y=1.465
+ $X2=0.39 $Y2=1.65
r103 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r104 31 35 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r105 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.975 $Y=1.765
+ $X2=2.975 $Y2=2.4
r106 24 30 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.565 $Y=1.65
+ $X2=2.475 $Y2=1.67
r107 23 25 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=2.885 $Y=1.65
+ $X2=2.975 $Y2=1.765
r108 23 24 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.885 $Y=1.65
+ $X2=2.565 $Y2=1.65
r109 20 30 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=2.475 $Y=1.765
+ $X2=2.475 $Y2=1.67
r110 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.475 $Y=1.765
+ $X2=2.475 $Y2=2.4
r111 19 29 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.115 $Y=1.65
+ $X2=2.025 $Y2=1.67
r112 18 30 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.385 $Y=1.65
+ $X2=2.475 $Y2=1.67
r113 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.385 $Y=1.65
+ $X2=2.115 $Y2=1.65
r114 15 29 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=2.025 $Y=1.765
+ $X2=2.025 $Y2=1.67
r115 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.025 $Y=1.765
+ $X2=2.025 $Y2=2.4
r116 14 28 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.665 $Y=1.65
+ $X2=1.575 $Y2=1.67
r117 13 29 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.935 $Y=1.65
+ $X2=2.025 $Y2=1.67
r118 13 14 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.935 $Y=1.65
+ $X2=1.665 $Y2=1.65
r119 10 28 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=1.575 $Y=1.765
+ $X2=1.575 $Y2=1.67
r120 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.575 $Y=1.765
+ $X2=1.575 $Y2=2.4
r121 9 36 31.3575 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.655 $Y=1.65
+ $X2=0.39 $Y2=1.65
r122 8 28 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.485 $Y=1.65
+ $X2=1.575 $Y2=1.67
r123 8 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.485 $Y=1.65
+ $X2=0.655 $Y2=1.65
r124 5 36 37.0701 $w=4.99e-07 $l=2.25278e-07 $layer=POLY_cond $X=0.565 $Y=1.765
+ $X2=0.39 $Y2=1.65
r125 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.565 $Y=1.765
+ $X2=0.565 $Y2=2.4
r126 1 34 41.8998 $w=4.99e-07 $l=2.11069e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.39 $Y2=1.465
r127 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 39
c87 1 0 4.66086e-20 $X=3.425 $Y=1.765
r88 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.88
+ $Y=1.385 $X2=4.88 $Y2=1.385
r89 39 41 9.04941 $w=5.06e-07 $l=9.5e-08 $layer=POLY_cond $X=4.785 $Y=1.492
+ $X2=4.88 $Y2=1.492
r90 38 39 0.952569 $w=5.06e-07 $l=1e-08 $layer=POLY_cond $X=4.775 $Y=1.492
+ $X2=4.785 $Y2=1.492
r91 37 38 40.0079 $w=5.06e-07 $l=4.2e-07 $layer=POLY_cond $X=4.355 $Y=1.492
+ $X2=4.775 $Y2=1.492
r92 36 37 2.85771 $w=5.06e-07 $l=3e-08 $layer=POLY_cond $X=4.325 $Y=1.492
+ $X2=4.355 $Y2=1.492
r93 34 36 11.9071 $w=5.06e-07 $l=1.25e-07 $layer=POLY_cond $X=4.2 $Y=1.492
+ $X2=4.325 $Y2=1.492
r94 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.2
+ $Y=1.385 $X2=4.2 $Y2=1.385
r95 32 34 27.1482 $w=5.06e-07 $l=2.85e-07 $layer=POLY_cond $X=3.915 $Y=1.492
+ $X2=4.2 $Y2=1.492
r96 31 32 3.81028 $w=5.06e-07 $l=4e-08 $layer=POLY_cond $X=3.875 $Y=1.492
+ $X2=3.915 $Y2=1.492
r97 30 31 37.1502 $w=5.06e-07 $l=3.9e-07 $layer=POLY_cond $X=3.485 $Y=1.492
+ $X2=3.875 $Y2=1.492
r98 29 30 5.71542 $w=5.06e-07 $l=6e-08 $layer=POLY_cond $X=3.425 $Y=1.492
+ $X2=3.485 $Y2=1.492
r99 26 42 4.98354 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.04 $Y=1.365
+ $X2=4.88 $Y2=1.365
r100 25 42 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.56 $Y=1.365
+ $X2=4.88 $Y2=1.365
r101 25 35 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.56 $Y=1.365
+ $X2=4.2 $Y2=1.365
r102 22 39 31.7097 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.785 $Y=1.22
+ $X2=4.785 $Y2=1.492
r103 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.785 $Y=1.22
+ $X2=4.785 $Y2=0.74
r104 19 38 31.7097 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.775 $Y=1.765
+ $X2=4.775 $Y2=1.492
r105 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.775 $Y=1.765
+ $X2=4.775 $Y2=2.4
r106 16 37 31.7097 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.355 $Y=1.22
+ $X2=4.355 $Y2=1.492
r107 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.355 $Y=1.22
+ $X2=4.355 $Y2=0.74
r108 13 36 31.7097 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.325 $Y=1.765
+ $X2=4.325 $Y2=1.492
r109 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.325 $Y=1.765
+ $X2=4.325 $Y2=2.4
r110 10 32 31.7097 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.915 $Y=1.22
+ $X2=3.915 $Y2=1.492
r111 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.915 $Y=1.22
+ $X2=3.915 $Y2=0.74
r112 7 31 31.7097 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.875 $Y2=1.492
r113 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.875 $Y2=2.4
r114 4 30 31.7097 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.485 $Y=1.22
+ $X2=3.485 $Y2=1.492
r115 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.485 $Y=1.22
+ $X2=3.485 $Y2=0.74
r116 1 29 31.7097 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.425 $Y=1.765
+ $X2=3.425 $Y2=1.492
r117 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.425 $Y=1.765
+ $X2=3.425 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_4%VPWR 1 2 3 10 12 18 24 28 30 35 45 46 52 55
r62 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r65 43 46 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r66 42 45 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r67 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 40 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=2.7 $Y2=3.33
r69 40 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 36 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.76 $Y2=3.33
r73 36 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 35 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=2.7 $Y2=3.33
r75 35 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 34 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 34 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r78 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 31 49 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r80 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 30 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=1.76 $Y2=3.33
r82 30 33 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 28 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r84 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r85 28 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 24 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.7 $Y=1.985 $X2=2.7
+ $Y2=2.815
r87 22 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=3.245 $X2=2.7
+ $Y2=3.33
r88 22 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.7 $Y=3.245 $X2=2.7
+ $Y2=2.815
r89 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.76 $Y=1.985
+ $X2=1.76 $Y2=2.815
r90 16 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=3.245
+ $X2=1.76 $Y2=3.33
r91 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.76 $Y=3.245
+ $X2=1.76 $Y2=2.815
r92 12 15 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.3 $Y=2.115 $X2=0.3
+ $Y2=2.815
r93 10 49 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.212 $Y2=3.33
r94 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.3 $Y=3.245 $X2=0.3
+ $Y2=2.815
r95 3 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.55
+ $Y=1.84 $X2=2.7 $Y2=2.815
r96 3 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.55
+ $Y=1.84 $X2=2.7 $Y2=1.985
r97 2 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.84 $X2=1.8 $Y2=2.815
r98 2 18 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.84 $X2=1.8 $Y2=1.985
r99 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.84 $X2=0.34 $Y2=2.815
r100 1 12 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.84 $X2=0.34 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_4%A_241_368# 1 2 3 4 5 18 22 23 26 30 35 38 39
+ 42 44 48 52 53
c96 39 0 9.04372e-20 $X=3.285 $Y=2.99
c97 35 0 2.55786e-19 $X=3.2 $Y=1.985
c98 26 0 1.20768e-19 $X=2.25 $Y=1.985
r99 48 51 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.04 $Y=1.985
+ $X2=5.04 $Y2=2.815
r100 46 51 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.04 $Y=2.905
+ $X2=5.04 $Y2=2.815
r101 45 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=2.99
+ $X2=4.1 $Y2=2.99
r102 44 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.915 $Y=2.99
+ $X2=5.04 $Y2=2.905
r103 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.915 $Y=2.99
+ $X2=4.185 $Y2=2.99
r104 40 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=2.905 $X2=4.1
+ $Y2=2.99
r105 40 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.1 $Y=2.905
+ $X2=4.1 $Y2=2.225
r106 38 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=2.99
+ $X2=4.1 $Y2=2.99
r107 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.015 $Y=2.99
+ $X2=3.285 $Y2=2.99
r108 35 37 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.16 $Y=1.985
+ $X2=3.16 $Y2=2.815
r109 33 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.16 $Y=2.905
+ $X2=3.285 $Y2=2.99
r110 33 37 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.16 $Y=2.905
+ $X2=3.16 $Y2=2.815
r111 32 35 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.16 $Y=1.65
+ $X2=3.16 $Y2=1.985
r112 31 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.335 $Y=1.565
+ $X2=2.21 $Y2=1.565
r113 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.035 $Y=1.565
+ $X2=3.16 $Y2=1.65
r114 30 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.035 $Y=1.565
+ $X2=2.335 $Y2=1.565
r115 26 28 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.21 $Y=1.985
+ $X2=2.21 $Y2=2.815
r116 24 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=1.65
+ $X2=2.21 $Y2=1.565
r117 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.21 $Y=1.65
+ $X2=2.21 $Y2=1.985
r118 22 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=1.565
+ $X2=2.21 $Y2=1.565
r119 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.085 $Y=1.565
+ $X2=1.435 $Y2=1.565
r120 18 20 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.31 $Y=1.985
+ $X2=1.31 $Y2=2.815
r121 16 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.31 $Y=1.65
+ $X2=1.435 $Y2=1.565
r122 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.31 $Y=1.65
+ $X2=1.31 $Y2=1.985
r123 5 51 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.85
+ $Y=1.84 $X2=5 $Y2=2.815
r124 5 48 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.85
+ $Y=1.84 $X2=5 $Y2=1.985
r125 4 42 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=3.95
+ $Y=1.84 $X2=4.1 $Y2=2.225
r126 3 37 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.05
+ $Y=1.84 $X2=3.2 $Y2=2.815
r127 3 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.05
+ $Y=1.84 $X2=3.2 $Y2=1.985
r128 2 28 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.84 $X2=2.25 $Y2=2.815
r129 2 26 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.84 $X2=2.25 $Y2=1.985
r130 1 20 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.84 $X2=1.35 $Y2=2.815
r131 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.84 $X2=1.35 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_4%Z 1 2 3 4 15 21 23 27 31 37 41 44
c51 44 0 1.82848e-19 $X=3.65 $Y=1.55
c52 41 0 1.40151e-19 $X=3.6 $Y=1.665
c53 21 0 4.66086e-20 $X=4.385 $Y=1.805
r54 41 46 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.65 $Y=1.665
+ $X2=3.65 $Y2=1.805
r55 41 44 5.79139 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.65 $Y=1.665
+ $X2=3.65 $Y2=1.55
r56 35 44 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=3.715 $Y=1.13
+ $X2=3.715 $Y2=1.55
r57 34 35 8.79174 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=3.74 $Y=0.95
+ $X2=3.74 $Y2=1.13
r58 31 34 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=3.74 $Y=0.89 $X2=3.74
+ $Y2=0.95
r59 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.55 $Y=1.97
+ $X2=4.55 $Y2=2.65
r60 25 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.55 $Y=1.89 $X2=4.55
+ $Y2=1.97
r61 24 31 0.964185 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=3.865 $Y=0.89
+ $X2=3.74 $Y2=0.89
r62 23 37 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.57 $Y=0.89 $X2=4.57
+ $Y2=0.8
r63 23 24 29.7714 $w=2.38e-07 $l=6.2e-07 $layer=LI1_cond $X=4.485 $Y=0.89
+ $X2=3.865 $Y2=0.89
r64 22 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=1.805
+ $X2=3.65 $Y2=1.805
r65 21 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.385 $Y=1.805
+ $X2=4.55 $Y2=1.89
r66 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.385 $Y=1.805
+ $X2=3.815 $Y2=1.805
r67 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.65 $Y=1.97
+ $X2=3.65 $Y2=2.65
r68 13 46 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=1.89
+ $X2=3.65 $Y2=1.805
r69 13 15 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.65 $Y=1.89 $X2=3.65
+ $Y2=1.97
r70 4 29 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.84 $X2=4.55 $Y2=2.65
r71 4 27 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.84 $X2=4.55 $Y2=1.97
r72 3 17 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.84 $X2=3.65 $Y2=2.65
r73 3 15 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.84 $X2=3.65 $Y2=1.97
r74 2 37 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.8
r75 1 34 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.37 $X2=3.7 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_4%VGND 1 2 3 10 12 16 20 23 24 26 27 28 44 45
c61 16 0 1.89802e-19 $X=1.98 $Y=0.515
r62 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r64 42 45 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r65 41 44 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r66 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r67 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r69 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r70 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r71 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r72 30 48 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r73 30 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r74 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r75 28 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r76 28 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r77 26 38 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.64
+ $Y2=0
r78 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.84
+ $Y2=0
r79 25 41 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=0 $X2=3.12
+ $Y2=0
r80 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0 $X2=2.84
+ $Y2=0
r81 23 35 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.68
+ $Y2=0
r82 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.98
+ $Y2=0
r83 22 38 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.64
+ $Y2=0
r84 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=1.98
+ $Y2=0
r85 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r86 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.515
r87 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r88 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.515
r89 10 48 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r90 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.515
r91 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.37 $X2=2.84 $Y2=0.515
r92 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.37 $X2=1.98 $Y2=0.515
r93 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_4%A_281_74# 1 2 3 4 5 18 20 21 24 26 28 29 30
+ 32 36 38 43
c82 38 0 1.72388e-19 $X=2.41 $Y=1.225
c83 21 0 3.63468e-19 $X=1.635 $Y=1.225
r84 42 43 8.64642 $w=3.43e-07 $l=1.7e-07 $layer=LI1_cond $X=4.135 $Y=0.427
+ $X2=4.305 $Y2=0.427
r85 34 36 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5 $Y=0.425 $X2=5
+ $Y2=0.68
r86 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.835 $Y=0.34
+ $X2=5 $Y2=0.425
r87 32 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.835 $Y=0.34
+ $X2=4.305 $Y2=0.34
r88 31 40 2.9551 $w=3.45e-07 $l=1.25e-07 $layer=LI1_cond $X=3.435 $Y=0.427
+ $X2=3.31 $Y2=0.427
r89 30 42 0.0668083 $w=3.43e-07 $l=2e-09 $layer=LI1_cond $X=4.133 $Y=0.427
+ $X2=4.135 $Y2=0.427
r90 30 31 23.3161 $w=3.43e-07 $l=6.98e-07 $layer=LI1_cond $X=4.133 $Y=0.427
+ $X2=3.435 $Y2=0.427
r91 28 40 4.08986 $w=2.5e-07 $l=1.73e-07 $layer=LI1_cond $X=3.31 $Y=0.6 $X2=3.31
+ $Y2=0.427
r92 28 29 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=3.31 $Y=0.6 $X2=3.31
+ $Y2=1.14
r93 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=1.225
+ $X2=2.41 $Y2=1.225
r94 26 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.185 $Y=1.225
+ $X2=3.31 $Y2=1.14
r95 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.185 $Y=1.225
+ $X2=2.495 $Y2=1.225
r96 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=1.14 $X2=2.41
+ $Y2=1.225
r97 22 24 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.41 $Y=1.14
+ $X2=2.41 $Y2=0.515
r98 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=1.225
+ $X2=2.41 $Y2=1.225
r99 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.325 $Y=1.225
+ $X2=1.635 $Y2=1.225
r100 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.55 $Y=1.14
+ $X2=1.635 $Y2=1.225
r101 16 18 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.55 $Y=1.14
+ $X2=1.55 $Y2=0.515
r102 5 36 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.68
r103 4 42 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.37 $X2=4.135 $Y2=0.515
r104 3 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.37 $X2=3.27 $Y2=0.515
r105 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.37 $X2=2.41 $Y2=0.515
r106 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.37 $X2=1.55 $Y2=0.515
.ends

