# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__nand3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.350000 1.095000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.820000 1.180000 7.075000 1.650000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.765000 1.350000 3.235000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.866500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685000 1.950000 5.850000 2.140000 ;
        RECT 3.750000 1.820000 5.850000 1.950000 ;
        RECT 4.130000 0.800000 5.345000 1.130000 ;
        RECT 4.925000 0.770000 5.345000 0.800000 ;
        RECT 4.925000 1.130000 5.155000 1.820000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.085000  0.580000 1.790000 0.670000 ;
      RECT 0.085000  0.670000 2.970000 0.750000 ;
      RECT 0.085000  0.750000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.785000 2.120000 ;
      RECT 0.115000  2.290000 0.445000 3.245000 ;
      RECT 0.425000  0.920000 0.755000 1.010000 ;
      RECT 0.425000  1.010000 3.770000 1.180000 ;
      RECT 0.615000  2.120000 0.785000 2.310000 ;
      RECT 0.615000  2.310000 6.230000 2.480000 ;
      RECT 0.935000  0.085000 1.280000 0.410000 ;
      RECT 0.955000  1.950000 1.435000 2.140000 ;
      RECT 1.265000  1.180000 1.435000 1.950000 ;
      RECT 1.460000  0.390000 1.790000 0.580000 ;
      RECT 1.460000  0.750000 2.970000 0.840000 ;
      RECT 1.490000  2.650000 2.565000 3.245000 ;
      RECT 1.970000  0.085000 2.460000 0.500000 ;
      RECT 2.640000  0.390000 2.970000 0.670000 ;
      RECT 3.135000  2.650000 3.630000 3.245000 ;
      RECT 3.140000  0.085000 3.470000 0.840000 ;
      RECT 3.600000  1.180000 3.770000 1.300000 ;
      RECT 3.600000  1.300000 4.610000 1.630000 ;
      RECT 3.700000  0.350000 7.565000 0.600000 ;
      RECT 3.700000  0.600000 4.030000 0.630000 ;
      RECT 4.580000  2.650000 5.400000 3.245000 ;
      RECT 5.515000  0.600000 7.565000 0.670000 ;
      RECT 5.945000  0.840000 7.415000 1.010000 ;
      RECT 5.970000  2.650000 7.565000 3.245000 ;
      RECT 6.060000  1.820000 7.415000 1.990000 ;
      RECT 6.060000  1.990000 6.230000 2.310000 ;
      RECT 6.400000  2.160000 7.565000 2.650000 ;
      RECT 7.245000  1.010000 7.415000 1.820000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__nand3b_4
END LIBRARY
