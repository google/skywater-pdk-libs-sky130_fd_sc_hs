* File: sky130_fd_sc_hs__dfrtp_4.pxi.spice
* Created: Thu Aug 27 20:38:53 2020
* 
x_PM_SKY130_FD_SC_HS__DFRTP_4%D N_D_c_280_n N_D_c_285_n N_D_c_286_n N_D_M1016_g
+ N_D_M1021_g D D D N_D_c_282_n N_D_c_283_n N_D_c_288_n
+ PM_SKY130_FD_SC_HS__DFRTP_4%D
x_PM_SKY130_FD_SC_HS__DFRTP_4%RESET_B N_RESET_B_M1009_g N_RESET_B_c_313_n
+ N_RESET_B_c_321_n N_RESET_B_c_322_n N_RESET_B_M1015_g N_RESET_B_c_314_n
+ N_RESET_B_M1034_g N_RESET_B_c_323_n N_RESET_B_c_324_n N_RESET_B_M1028_g
+ N_RESET_B_c_315_n N_RESET_B_c_326_n N_RESET_B_M1002_g N_RESET_B_M1031_g
+ N_RESET_B_c_317_n N_RESET_B_c_328_n N_RESET_B_c_329_n N_RESET_B_c_330_n
+ N_RESET_B_c_331_n N_RESET_B_c_332_n N_RESET_B_c_333_n N_RESET_B_c_334_n
+ N_RESET_B_c_335_n RESET_B N_RESET_B_c_336_n N_RESET_B_c_318_n
+ N_RESET_B_c_319_n N_RESET_B_c_338_n PM_SKY130_FD_SC_HS__DFRTP_4%RESET_B
x_PM_SKY130_FD_SC_HS__DFRTP_4%CLK N_CLK_M1026_g N_CLK_c_527_n N_CLK_M1004_g CLK
+ PM_SKY130_FD_SC_HS__DFRTP_4%CLK
x_PM_SKY130_FD_SC_HS__DFRTP_4%A_494_366# N_A_494_366#_M1012_d
+ N_A_494_366#_M1010_d N_A_494_366#_c_589_n N_A_494_366#_c_590_n
+ N_A_494_366#_M1027_g N_A_494_366#_c_570_n N_A_494_366#_c_571_n
+ N_A_494_366#_M1035_g N_A_494_366#_c_573_n N_A_494_366#_M1006_g
+ N_A_494_366#_c_574_n N_A_494_366#_c_575_n N_A_494_366#_c_593_n
+ N_A_494_366#_M1020_g N_A_494_366#_c_576_n N_A_494_366#_c_577_n
+ N_A_494_366#_c_595_n N_A_494_366#_c_596_n N_A_494_366#_c_578_n
+ N_A_494_366#_c_579_n N_A_494_366#_c_580_n N_A_494_366#_c_581_n
+ N_A_494_366#_c_582_n N_A_494_366#_c_583_n N_A_494_366#_c_584_n
+ N_A_494_366#_c_585_n N_A_494_366#_c_586_n N_A_494_366#_c_587_n
+ N_A_494_366#_c_588_n PM_SKY130_FD_SC_HS__DFRTP_4%A_494_366#
x_PM_SKY130_FD_SC_HS__DFRTP_4%A_834_355# N_A_834_355#_M1017_d
+ N_A_834_355#_M1005_d N_A_834_355#_c_774_n N_A_834_355#_M1019_g
+ N_A_834_355#_M1025_g N_A_834_355#_c_772_n N_A_834_355#_c_807_n
+ N_A_834_355#_c_773_n N_A_834_355#_c_809_n N_A_834_355#_c_817_p
+ N_A_834_355#_c_793_n N_A_834_355#_c_778_n
+ PM_SKY130_FD_SC_HS__DFRTP_4%A_834_355#
x_PM_SKY130_FD_SC_HS__DFRTP_4%A_313_74# N_A_313_74#_M1026_s N_A_313_74#_M1004_s
+ N_A_313_74#_c_874_n N_A_313_74#_M1010_g N_A_313_74#_c_859_n
+ N_A_313_74#_M1012_g N_A_313_74#_c_860_n N_A_313_74#_c_875_n
+ N_A_313_74#_c_876_n N_A_313_74#_c_877_n N_A_313_74#_c_861_n
+ N_A_313_74#_M1001_g N_A_313_74#_c_878_n N_A_313_74#_c_879_n
+ N_A_313_74#_c_880_n N_A_313_74#_M1029_g N_A_313_74#_c_881_n
+ N_A_313_74#_c_882_n N_A_313_74#_c_862_n N_A_313_74#_M1011_g
+ N_A_313_74#_c_863_n N_A_313_74#_M1037_g N_A_313_74#_c_865_n
+ N_A_313_74#_c_866_n N_A_313_74#_c_886_n N_A_313_74#_c_867_n
+ N_A_313_74#_c_868_n N_A_313_74#_c_869_n N_A_313_74#_c_870_n
+ N_A_313_74#_c_871_n N_A_313_74#_c_888_n N_A_313_74#_c_889_n
+ N_A_313_74#_c_872_n N_A_313_74#_c_890_n N_A_313_74#_c_891_n
+ N_A_313_74#_c_892_n N_A_313_74#_c_873_n PM_SKY130_FD_SC_HS__DFRTP_4%A_313_74#
x_PM_SKY130_FD_SC_HS__DFRTP_4%A_699_463# N_A_699_463#_M1001_d
+ N_A_699_463#_M1027_d N_A_699_463#_M1028_d N_A_699_463#_c_1086_n
+ N_A_699_463#_M1017_g N_A_699_463#_c_1095_n N_A_699_463#_M1005_g
+ N_A_699_463#_c_1087_n N_A_699_463#_c_1088_n N_A_699_463#_c_1089_n
+ N_A_699_463#_c_1090_n N_A_699_463#_c_1110_n N_A_699_463#_c_1098_n
+ N_A_699_463#_c_1091_n N_A_699_463#_c_1092_n N_A_699_463#_c_1093_n
+ N_A_699_463#_c_1094_n N_A_699_463#_c_1100_n
+ PM_SKY130_FD_SC_HS__DFRTP_4%A_699_463#
x_PM_SKY130_FD_SC_HS__DFRTP_4%A_1678_395# N_A_1678_395#_M1032_d
+ N_A_1678_395#_M1002_d N_A_1678_395#_c_1227_n N_A_1678_395#_c_1228_n
+ N_A_1678_395#_M1000_g N_A_1678_395#_M1023_g N_A_1678_395#_c_1220_n
+ N_A_1678_395#_c_1230_n N_A_1678_395#_c_1221_n N_A_1678_395#_c_1231_n
+ N_A_1678_395#_c_1232_n N_A_1678_395#_c_1233_n N_A_1678_395#_c_1222_n
+ N_A_1678_395#_c_1223_n N_A_1678_395#_c_1224_n N_A_1678_395#_c_1225_n
+ N_A_1678_395#_c_1235_n N_A_1678_395#_c_1226_n
+ PM_SKY130_FD_SC_HS__DFRTP_4%A_1678_395#
x_PM_SKY130_FD_SC_HS__DFRTP_4%A_1350_392# N_A_1350_392#_M1006_d
+ N_A_1350_392#_M1011_d N_A_1350_392#_M1032_g N_A_1350_392#_c_1357_n
+ N_A_1350_392#_c_1358_n N_A_1350_392#_M1008_g N_A_1350_392#_c_1344_n
+ N_A_1350_392#_c_1360_n N_A_1350_392#_c_1361_n N_A_1350_392#_M1018_g
+ N_A_1350_392#_c_1345_n N_A_1350_392#_c_1363_n N_A_1350_392#_c_1364_n
+ N_A_1350_392#_M1030_g N_A_1350_392#_c_1346_n N_A_1350_392#_M1022_g
+ N_A_1350_392#_c_1347_n N_A_1350_392#_c_1348_n N_A_1350_392#_c_1349_n
+ N_A_1350_392#_c_1350_n N_A_1350_392#_c_1393_n N_A_1350_392#_c_1351_n
+ N_A_1350_392#_c_1352_n N_A_1350_392#_c_1380_n N_A_1350_392#_c_1368_n
+ N_A_1350_392#_c_1353_n N_A_1350_392#_c_1354_n N_A_1350_392#_c_1355_n
+ N_A_1350_392#_c_1356_n PM_SKY130_FD_SC_HS__DFRTP_4%A_1350_392#
x_PM_SKY130_FD_SC_HS__DFRTP_4%A_2010_409# N_A_2010_409#_M1022_d
+ N_A_2010_409#_M1018_d N_A_2010_409#_c_1523_n N_A_2010_409#_M1007_g
+ N_A_2010_409#_c_1509_n N_A_2010_409#_c_1524_n N_A_2010_409#_M1013_g
+ N_A_2010_409#_M1003_g N_A_2010_409#_c_1511_n N_A_2010_409#_c_1512_n
+ N_A_2010_409#_M1024_g N_A_2010_409#_c_1526_n N_A_2010_409#_M1014_g
+ N_A_2010_409#_M1033_g N_A_2010_409#_c_1527_n N_A_2010_409#_M1036_g
+ N_A_2010_409#_M1038_g N_A_2010_409#_c_1516_n N_A_2010_409#_c_1529_n
+ N_A_2010_409#_c_1517_n N_A_2010_409#_c_1518_n N_A_2010_409#_c_1519_n
+ N_A_2010_409#_c_1520_n N_A_2010_409#_c_1521_n N_A_2010_409#_c_1522_n
+ PM_SKY130_FD_SC_HS__DFRTP_4%A_2010_409#
x_PM_SKY130_FD_SC_HS__DFRTP_4%VPWR N_VPWR_M1016_s N_VPWR_M1015_d N_VPWR_M1004_d
+ N_VPWR_M1019_d N_VPWR_M1005_s N_VPWR_M1000_d N_VPWR_M1008_d N_VPWR_M1030_s
+ N_VPWR_M1013_s N_VPWR_M1036_s N_VPWR_c_1641_n N_VPWR_c_1642_n N_VPWR_c_1643_n
+ N_VPWR_c_1644_n N_VPWR_c_1645_n N_VPWR_c_1646_n N_VPWR_c_1647_n
+ N_VPWR_c_1648_n N_VPWR_c_1649_n N_VPWR_c_1650_n N_VPWR_c_1651_n
+ N_VPWR_c_1652_n N_VPWR_c_1653_n N_VPWR_c_1654_n N_VPWR_c_1655_n
+ N_VPWR_c_1656_n N_VPWR_c_1657_n N_VPWR_c_1658_n VPWR N_VPWR_c_1659_n
+ N_VPWR_c_1660_n N_VPWR_c_1661_n N_VPWR_c_1662_n N_VPWR_c_1663_n
+ N_VPWR_c_1664_n N_VPWR_c_1665_n N_VPWR_c_1666_n N_VPWR_c_1667_n
+ N_VPWR_c_1668_n N_VPWR_c_1669_n N_VPWR_c_1640_n
+ PM_SKY130_FD_SC_HS__DFRTP_4%VPWR
x_PM_SKY130_FD_SC_HS__DFRTP_4%A_37_78# N_A_37_78#_M1021_s N_A_37_78#_M1001_s
+ N_A_37_78#_M1016_d N_A_37_78#_M1027_s N_A_37_78#_c_1805_n N_A_37_78#_c_1806_n
+ N_A_37_78#_c_1813_n N_A_37_78#_c_1807_n N_A_37_78#_c_1814_n
+ N_A_37_78#_c_1808_n N_A_37_78#_c_1809_n N_A_37_78#_c_1810_n
+ N_A_37_78#_c_1811_n N_A_37_78#_c_1816_n N_A_37_78#_c_1817_n
+ N_A_37_78#_c_1818_n N_A_37_78#_c_1819_n PM_SKY130_FD_SC_HS__DFRTP_4%A_37_78#
x_PM_SKY130_FD_SC_HS__DFRTP_4%Q N_Q_M1003_s N_Q_M1033_s N_Q_M1007_d N_Q_M1014_d
+ N_Q_c_1939_n N_Q_c_1940_n N_Q_c_1941_n N_Q_c_1932_n N_Q_c_1933_n N_Q_c_1934_n
+ N_Q_c_1942_n N_Q_c_1935_n N_Q_c_1936_n N_Q_c_1937_n Q
+ PM_SKY130_FD_SC_HS__DFRTP_4%Q
x_PM_SKY130_FD_SC_HS__DFRTP_4%VGND N_VGND_M1009_d N_VGND_M1026_d N_VGND_M1034_d
+ N_VGND_M1023_d N_VGND_M1022_s N_VGND_M1003_d N_VGND_M1024_d N_VGND_M1038_d
+ N_VGND_c_2006_n N_VGND_c_2007_n N_VGND_c_2008_n N_VGND_c_2009_n
+ N_VGND_c_2010_n N_VGND_c_2011_n N_VGND_c_2012_n N_VGND_c_2013_n
+ N_VGND_c_2014_n N_VGND_c_2015_n N_VGND_c_2016_n N_VGND_c_2017_n VGND
+ N_VGND_c_2018_n N_VGND_c_2019_n N_VGND_c_2020_n N_VGND_c_2021_n
+ N_VGND_c_2022_n N_VGND_c_2023_n N_VGND_c_2024_n N_VGND_c_2025_n
+ N_VGND_c_2026_n N_VGND_c_2027_n N_VGND_c_2028_n N_VGND_c_2029_n
+ PM_SKY130_FD_SC_HS__DFRTP_4%VGND
cc_1 VNB N_D_c_280_n 0.0407866f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.81
cc_2 VNB N_D_M1021_g 0.0286444f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_3 VNB N_D_c_282_n 0.0249067f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_283_n 0.0295836f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB N_RESET_B_M1009_g 0.0302022f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.01
cc_6 VNB N_RESET_B_c_313_n 0.0274408f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_7 VNB N_RESET_B_c_314_n 0.0174763f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_RESET_B_c_315_n 0.021059f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1
cc_9 VNB N_RESET_B_M1031_g 0.0519609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_RESET_B_c_317_n 0.0175891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_RESET_B_c_318_n 0.0317115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_RESET_B_c_319_n 0.00562946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_CLK_M1026_g 0.0265896f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.01
cc_14 VNB N_CLK_c_527_n 0.0328676f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_15 VNB CLK 0.00638992f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1
cc_16 VNB N_A_494_366#_c_570_n 0.00917687f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A_494_366#_c_571_n 0.021321f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_18 VNB N_A_494_366#_M1035_g 0.0241841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_494_366#_c_573_n 0.0216455f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.165
cc_20 VNB N_A_494_366#_c_574_n 0.0206494f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1
cc_21 VNB N_A_494_366#_c_575_n 0.00999606f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.845
cc_22 VNB N_A_494_366#_c_576_n 0.0103565f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_23 VNB N_A_494_366#_c_577_n 0.0395914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_494_366#_c_578_n 0.00519588f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_25 VNB N_A_494_366#_c_579_n 0.0255302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_494_366#_c_580_n 0.00585827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_494_366#_c_581_n 0.00192671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_494_366#_c_582_n 0.0117871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_494_366#_c_583_n 0.00162301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_494_366#_c_584_n 0.0109807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_494_366#_c_585_n 0.0026267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_494_366#_c_586_n 0.030848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_494_366#_c_587_n 0.00738738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_494_366#_c_588_n 0.00971843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_834_355#_M1025_g 0.0367823f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VNB N_A_834_355#_c_772_n 0.00382242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_834_355#_c_773_n 0.00906432f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.845
cc_38 VNB N_A_313_74#_c_859_n 0.0212781f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_39 VNB N_A_313_74#_c_860_n 0.0483384f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_40 VNB N_A_313_74#_c_861_n 0.017907f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_41 VNB N_A_313_74#_c_862_n 0.0368495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_313_74#_c_863_n 0.0331371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_313_74#_M1037_g 0.0499146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_313_74#_c_865_n 0.0144643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_313_74#_c_866_n 0.00954314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_313_74#_c_867_n 0.011229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_313_74#_c_868_n 0.00958559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_313_74#_c_869_n 0.0046226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_313_74#_c_870_n 5.44847e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_313_74#_c_871_n 0.016061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_313_74#_c_872_n 0.00536974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_313_74#_c_873_n 0.00625184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_699_463#_c_1086_n 0.0239206f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_54 VNB N_A_699_463#_c_1087_n 0.0175129f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.165
cc_55 VNB N_A_699_463#_c_1088_n 0.0496697f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_56 VNB N_A_699_463#_c_1089_n 0.00824647f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_57 VNB N_A_699_463#_c_1090_n 0.00401724f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=1.845
cc_58 VNB N_A_699_463#_c_1091_n 0.00102843f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.165
cc_59 VNB N_A_699_463#_c_1092_n 0.00109066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_699_463#_c_1093_n 0.0134696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_699_463#_c_1094_n 0.00277203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1678_395#_M1023_g 0.0226108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1678_395#_c_1220_n 0.0147871f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=1.165
cc_64 VNB N_A_1678_395#_c_1221_n 0.0161902f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_65 VNB N_A_1678_395#_c_1222_n 0.0100185f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.295
cc_66 VNB N_A_1678_395#_c_1223_n 0.00724983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1678_395#_c_1224_n 0.00408177f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.845
cc_68 VNB N_A_1678_395#_c_1225_n 0.0315912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1678_395#_c_1226_n 0.00985953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1350_392#_M1032_g 0.0443312f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_71 VNB N_A_1350_392#_c_1344_n 0.00790233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1350_392#_c_1345_n 0.0119253f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_73 VNB N_A_1350_392#_c_1346_n 0.0144823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1350_392#_c_1347_n 0.0103327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1350_392#_c_1348_n 0.00465184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1350_392#_c_1349_n 0.0189463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1350_392#_c_1350_n 0.0167302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1350_392#_c_1351_n 0.00538628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1350_392#_c_1352_n 0.0041539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1350_392#_c_1353_n 0.00737056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1350_392#_c_1354_n 0.00664015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1350_392#_c_1355_n 0.00100027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1350_392#_c_1356_n 0.0239677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2010_409#_c_1509_n 0.0142504f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_85 VNB N_A_2010_409#_M1003_g 0.0250105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2010_409#_c_1511_n 0.0271444f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_87 VNB N_A_2010_409#_c_1512_n 0.028357f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_88 VNB N_A_2010_409#_M1024_g 0.0223949f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_89 VNB N_A_2010_409#_M1033_g 0.02888f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_90 VNB N_A_2010_409#_M1038_g 0.0378399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2010_409#_c_1516_n 0.0119979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2010_409#_c_1517_n 0.00142943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2010_409#_c_1518_n 0.00371217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2010_409#_c_1519_n 0.0128657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2010_409#_c_1520_n 0.0109985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2010_409#_c_1521_n 0.0048999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2010_409#_c_1522_n 0.0647225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VPWR_c_1640_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_37_78#_c_1805_n 0.00234939f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_100 VNB N_A_37_78#_c_1806_n 0.0151278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_37_78#_c_1807_n 0.0027805f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_102 VNB N_A_37_78#_c_1808_n 0.00608807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_37_78#_c_1809_n 0.00178054f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_104 VNB N_A_37_78#_c_1810_n 0.00406071f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_105 VNB N_A_37_78#_c_1811_n 0.0222792f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_106 VNB N_Q_c_1932_n 0.00250883f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1
cc_107 VNB N_Q_c_1933_n 0.00280896f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_108 VNB N_Q_c_1934_n 0.00323677f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.01
cc_109 VNB N_Q_c_1935_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_Q_c_1936_n 0.00131414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_Q_c_1937_n 2.04518e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB Q 0.0222191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2006_n 0.0112006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2007_n 0.00961509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2008_n 0.0151521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2009_n 0.0133586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2010_n 0.0179738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2011_n 0.00503034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2012_n 0.0117082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2013_n 0.0382127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2014_n 0.0320339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2015_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2016_n 0.0344576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2017_n 0.00528956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2018_n 0.0224468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2019_n 0.0622418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2020_n 0.0798951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2021_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2022_n 0.0187248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2023_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2024_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2025_n 0.0162053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2026_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2027_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2028_n 0.00606636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2029_n 0.747947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VPB N_D_c_280_n 0.0132401f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.81
cc_138 VPB N_D_c_285_n 0.0381729f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.245
cc_139 VPB N_D_c_286_n 0.0179054f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.465
cc_140 VPB N_D_c_283_n 0.0247385f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_141 VPB N_D_c_288_n 0.0231943f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_142 VPB N_RESET_B_c_313_n 0.0234263f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_143 VPB N_RESET_B_c_321_n 0.0179997f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_144 VPB N_RESET_B_c_322_n 0.0236024f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.6
cc_145 VPB N_RESET_B_c_323_n 0.0095874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_RESET_B_c_324_n 0.0223373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_c_315_n 7.13987e-19 $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1
cc_148 VPB N_RESET_B_c_326_n 0.0521136f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.845
cc_149 VPB N_RESET_B_M1031_g 0.0152075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_328_n 0.0106508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_329_n 0.0230319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_330_n 0.00380423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_331_n 0.0267148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_RESET_B_c_332_n 0.00376976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_RESET_B_c_333_n 0.0151408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_RESET_B_c_334_n 0.00293589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_RESET_B_c_335_n 0.00604009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_RESET_B_c_336_n 0.0469968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_RESET_B_c_319_n 9.23273e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_c_338_n 0.0286678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_CLK_c_527_n 0.0239557f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.465
cc_162 VPB CLK 0.00474195f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_163 VPB N_A_494_366#_c_589_n 0.0160416f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_164 VPB N_A_494_366#_c_590_n 0.01982f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.6
cc_165 VPB N_A_494_366#_c_570_n 0.00974149f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_166 VPB N_A_494_366#_c_571_n 0.00693897f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_167 VPB N_A_494_366#_c_593_n 0.0671551f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_168 VPB N_A_494_366#_c_576_n 2.57762e-19 $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_169 VPB N_A_494_366#_c_595_n 0.00324726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_494_366#_c_596_n 0.00105171f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_171 VPB N_A_494_366#_c_580_n 0.00688356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_494_366#_c_583_n 0.00100773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_494_366#_c_588_n 0.0191897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_834_355#_c_774_n 0.0687453f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_175 VPB N_A_834_355#_M1025_g 0.00601276f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_176 VPB N_A_834_355#_c_772_n 0.00190944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_834_355#_c_773_n 0.00257559f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.845
cc_178 VPB N_A_834_355#_c_778_n 0.00722631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_313_74#_c_874_n 0.0143065f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_180 VPB N_A_313_74#_c_875_n 0.0769393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_313_74#_c_876_n 0.0552222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_313_74#_c_877_n 0.0125211f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.165
cc_183 VPB N_A_313_74#_c_878_n 0.00711171f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.845
cc_184 VPB N_A_313_74#_c_879_n 0.01637f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_185 VPB N_A_313_74#_c_880_n 0.0143055f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_186 VPB N_A_313_74#_c_881_n 0.107363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_313_74#_c_882_n 0.0379082f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_188 VPB N_A_313_74#_c_862_n 0.0348925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_313_74#_c_863_n 0.0503144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_313_74#_c_866_n 0.0205253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_313_74#_c_886_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_313_74#_c_868_n 0.00365578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_313_74#_c_888_n 0.00410718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_313_74#_c_889_n 0.004254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_313_74#_c_890_n 0.00727491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_313_74#_c_891_n 0.00400849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_313_74#_c_892_n 0.0467154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_699_463#_c_1095_n 0.0286139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_699_463#_c_1089_n 0.00436657f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_200 VPB N_A_699_463#_c_1090_n 0.0109849f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.845
cc_201 VPB N_A_699_463#_c_1098_n 0.00239748f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.845
cc_202 VPB N_A_699_463#_c_1091_n 0.00424035f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.165
cc_203 VPB N_A_699_463#_c_1100_n 0.00353943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1678_395#_c_1227_n 0.00843909f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_205 VPB N_A_1678_395#_c_1228_n 0.0213158f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.6
cc_206 VPB N_A_1678_395#_c_1220_n 0.017829f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.165
cc_207 VPB N_A_1678_395#_c_1230_n 0.00940749f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_208 VPB N_A_1678_395#_c_1231_n 0.00319167f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.845
cc_209 VPB N_A_1678_395#_c_1232_n 0.00693697f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.845
cc_210 VPB N_A_1678_395#_c_1233_n 0.00169772f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=2.01
cc_211 VPB N_A_1678_395#_c_1223_n 0.00167634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1678_395#_c_1235_n 0.0100342f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1350_392#_c_1357_n 0.0301229f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_214 VPB N_A_1350_392#_c_1358_n 0.0208013f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_215 VPB N_A_1350_392#_c_1344_n 0.00374484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1350_392#_c_1360_n 0.00873449f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_217 VPB N_A_1350_392#_c_1361_n 0.0205027f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_218 VPB N_A_1350_392#_c_1345_n 0.00385745f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.845
cc_219 VPB N_A_1350_392#_c_1363_n 0.00915965f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.165
cc_220 VPB N_A_1350_392#_c_1364_n 0.0210658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1350_392#_c_1347_n 8.59645e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1350_392#_c_1348_n 0.00184123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1350_392#_c_1351_n 0.0164504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1350_392#_c_1368_n 0.00772571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1350_392#_c_1353_n 0.00974213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1350_392#_c_1354_n 2.91644e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1350_392#_c_1355_n 3.14732e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1350_392#_c_1356_n 0.00359861f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_2010_409#_c_1523_n 0.0168955f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_230 VPB N_A_2010_409#_c_1524_n 0.0176613f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_231 VPB N_A_2010_409#_c_1512_n 0.00975576f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_232 VPB N_A_2010_409#_c_1526_n 0.017171f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=2.01
cc_233 VPB N_A_2010_409#_c_1527_n 0.017675f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_234 VPB N_A_2010_409#_c_1516_n 0.00731318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_2010_409#_c_1529_n 0.00457997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_2010_409#_c_1522_n 0.0163813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1641_n 0.0104926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1642_n 0.0319294f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.035
cc_239 VPB N_VPWR_c_1643_n 0.012732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1644_n 0.0036638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1645_n 0.00946291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1646_n 0.00703496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1647_n 0.0199844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1648_n 0.0124761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1649_n 0.00722026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1650_n 0.0122465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1651_n 0.0149023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1652_n 0.0511093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1653_n 0.0667644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1654_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1655_n 0.020793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1656_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1657_n 0.0184712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1658_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1659_n 0.0205885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1660_n 0.0210058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1661_n 0.0595607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1662_n 0.0303917f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1663_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1664_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1665_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1666_n 0.00613849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1667_n 0.00436844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1668_n 0.00623693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1669_n 0.0135346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1640_n 0.139332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_37_78#_c_1806_n 0.0108264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_37_78#_c_1813_n 0.00346984f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_269 VPB N_A_37_78#_c_1814_n 0.00624613f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=2.01
cc_270 VPB N_A_37_78#_c_1810_n 0.0051551f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_271 VPB N_A_37_78#_c_1816_n 0.00798703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_37_78#_c_1817_n 0.0112223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_37_78#_c_1818_n 0.00255485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_37_78#_c_1819_n 0.00924367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_Q_c_1939_n 0.00289698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_Q_c_1940_n 0.00522595f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_277 VPB N_Q_c_1941_n 0.00246435f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_278 VPB N_Q_c_1942_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB Q 0.0128167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 N_D_M1021_g N_RESET_B_M1009_g 0.0204989f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_281 N_D_c_280_n N_RESET_B_c_313_n 0.0204989f $X=0.42 $Y=1.81 $X2=0 $Y2=0
cc_282 N_D_c_285_n N_RESET_B_c_321_n 0.0253834f $X=0.515 $Y=2.245 $X2=0 $Y2=0
cc_283 N_D_c_286_n N_RESET_B_c_322_n 0.00917787f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_284 N_D_c_282_n N_RESET_B_c_318_n 0.0204989f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_285 N_D_c_288_n N_RESET_B_c_338_n 0.0204989f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_286 N_D_c_286_n N_VPWR_c_1642_n 0.00729224f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_287 N_D_c_283_n N_VPWR_c_1642_n 0.0134569f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_288 N_D_c_288_n N_VPWR_c_1642_n 7.3436e-19 $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_289 N_D_c_286_n N_VPWR_c_1659_n 0.00444469f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_290 N_D_c_285_n N_VPWR_c_1640_n 3.7828e-19 $X=0.515 $Y=2.245 $X2=0 $Y2=0
cc_291 N_D_c_286_n N_VPWR_c_1640_n 0.00857482f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_292 N_D_M1021_g N_A_37_78#_c_1805_n 0.0116103f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_293 N_D_c_283_n N_A_37_78#_c_1805_n 0.00144733f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_294 N_D_M1021_g N_A_37_78#_c_1806_n 0.0152984f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_295 N_D_c_283_n N_A_37_78#_c_1806_n 0.0891656f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_296 N_D_M1021_g N_A_37_78#_c_1811_n 0.00807807f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_297 N_D_c_282_n N_A_37_78#_c_1811_n 0.00188146f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_298 N_D_c_283_n N_A_37_78#_c_1811_n 0.0285087f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_299 N_D_c_285_n N_A_37_78#_c_1816_n 0.00687401f $X=0.515 $Y=2.245 $X2=0 $Y2=0
cc_300 N_D_c_286_n N_A_37_78#_c_1816_n 0.00810441f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_301 N_D_M1021_g N_VGND_c_2014_n 0.00429844f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_302 N_D_M1021_g N_VGND_c_2029_n 0.00539454f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_303 N_RESET_B_c_318_n N_CLK_M1026_g 0.0027096f $X=1.155 $Y=1.295 $X2=0 $Y2=0
cc_304 N_RESET_B_c_313_n N_CLK_c_527_n 0.00594633f $X=1.09 $Y=1.91 $X2=0 $Y2=0
cc_305 N_RESET_B_c_329_n N_CLK_c_527_n 0.0054633f $X=5.375 $Y=2.035 $X2=0 $Y2=0
cc_306 N_RESET_B_c_318_n N_CLK_c_527_n 0.00678299f $X=1.155 $Y=1.295 $X2=0 $Y2=0
cc_307 N_RESET_B_c_329_n CLK 0.0159129f $X=5.375 $Y=2.035 $X2=0 $Y2=0
cc_308 N_RESET_B_c_329_n N_A_494_366#_c_589_n 0.00345345f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_309 N_RESET_B_c_329_n N_A_494_366#_c_570_n 0.00443957f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_310 N_RESET_B_c_329_n N_A_494_366#_c_571_n 3.82592e-19 $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_311 N_RESET_B_c_331_n N_A_494_366#_c_593_n 0.0037737f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_312 N_RESET_B_c_329_n N_A_494_366#_c_595_n 0.0049998f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_313 N_RESET_B_c_329_n N_A_494_366#_c_596_n 0.0295434f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_314 N_RESET_B_c_314_n N_A_494_366#_c_578_n 0.0108891f $X=4.765 $Y=1.185 $X2=0
+ $Y2=0
cc_315 N_RESET_B_c_331_n N_A_494_366#_c_580_n 0.0224618f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_316 N_RESET_B_c_329_n N_A_494_366#_c_583_n 0.00693564f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_317 N_RESET_B_c_314_n N_A_494_366#_c_585_n 3.16315e-19 $X=4.765 $Y=1.185
+ $X2=0 $Y2=0
cc_318 N_RESET_B_c_329_n N_A_494_366#_c_588_n 2.80857e-19 $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_319 N_RESET_B_c_323_n N_A_834_355#_c_774_n 0.00319024f $X=4.87 $Y=2.15 $X2=0
+ $Y2=0
cc_320 N_RESET_B_c_324_n N_A_834_355#_c_774_n 0.0138579f $X=4.87 $Y=2.24 $X2=0
+ $Y2=0
cc_321 N_RESET_B_c_328_n N_A_834_355#_c_774_n 0.0215869f $X=4.87 $Y=1.835 $X2=0
+ $Y2=0
cc_322 N_RESET_B_c_329_n N_A_834_355#_c_774_n 0.00908008f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_323 N_RESET_B_c_314_n N_A_834_355#_M1025_g 0.0417267f $X=4.765 $Y=1.185 $X2=0
+ $Y2=0
cc_324 N_RESET_B_c_315_n N_A_834_355#_M1025_g 0.0107658f $X=4.885 $Y=1.67 $X2=0
+ $Y2=0
cc_325 N_RESET_B_c_328_n N_A_834_355#_M1025_g 0.00382675f $X=4.87 $Y=1.835 $X2=0
+ $Y2=0
cc_326 N_RESET_B_c_314_n N_A_834_355#_c_772_n 0.00472366f $X=4.765 $Y=1.185
+ $X2=0 $Y2=0
cc_327 N_RESET_B_c_315_n N_A_834_355#_c_772_n 0.00104148f $X=4.885 $Y=1.67 $X2=0
+ $Y2=0
cc_328 N_RESET_B_c_328_n N_A_834_355#_c_772_n 8.0459e-19 $X=4.87 $Y=1.835 $X2=0
+ $Y2=0
cc_329 N_RESET_B_c_329_n N_A_834_355#_c_772_n 0.0222661f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_330 N_RESET_B_c_331_n N_A_834_355#_c_773_n 0.00270439f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_331 N_RESET_B_c_332_n N_A_834_355#_c_773_n 4.50751e-19 $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_332 N_RESET_B_c_333_n N_A_834_355#_c_773_n 0.00890751f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_333 N_RESET_B_c_314_n N_A_834_355#_c_793_n 0.0136619f $X=4.765 $Y=1.185 $X2=0
+ $Y2=0
cc_334 N_RESET_B_c_317_n N_A_834_355#_c_793_n 0.00316016f $X=4.885 $Y=1.26 $X2=0
+ $Y2=0
cc_335 N_RESET_B_c_331_n N_A_834_355#_c_778_n 0.0278833f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_336 N_RESET_B_c_332_n N_A_834_355#_c_778_n 0.0020002f $X=5.665 $Y=2.035 $X2=0
+ $Y2=0
cc_337 N_RESET_B_c_333_n N_A_834_355#_c_778_n 0.00333678f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_338 N_RESET_B_c_329_n N_A_313_74#_M1004_s 0.00115255f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_339 N_RESET_B_c_329_n N_A_313_74#_c_874_n 0.00773946f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_340 N_RESET_B_c_329_n N_A_313_74#_c_875_n 0.00334754f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_341 N_RESET_B_c_329_n N_A_313_74#_c_880_n 0.00253485f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_342 N_RESET_B_c_324_n N_A_313_74#_c_881_n 0.00990349f $X=4.87 $Y=2.24 $X2=0
+ $Y2=0
cc_343 N_RESET_B_c_331_n N_A_313_74#_c_862_n 0.0221149f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_344 N_RESET_B_c_329_n N_A_313_74#_c_866_n 3.88441e-19 $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_345 N_RESET_B_M1009_g N_A_313_74#_c_867_n 0.00344772f $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_346 N_RESET_B_c_329_n N_A_313_74#_c_868_n 8.85602e-19 $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_347 N_RESET_B_c_318_n N_A_313_74#_c_868_n 0.00656198f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_348 N_RESET_B_c_319_n N_A_313_74#_c_868_n 0.049377f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_349 N_RESET_B_c_329_n N_A_313_74#_c_870_n 0.00130818f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_350 N_RESET_B_c_331_n N_A_313_74#_c_888_n 0.0254407f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_351 N_RESET_B_c_331_n N_A_313_74#_c_889_n 0.0163819f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_352 N_RESET_B_M1009_g N_A_313_74#_c_872_n 0.00291406f $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_353 N_RESET_B_c_319_n N_A_313_74#_c_872_n 8.29766e-19 $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_354 N_RESET_B_c_313_n N_A_313_74#_c_890_n 0.00299847f $X=1.09 $Y=1.91 $X2=0
+ $Y2=0
cc_355 N_RESET_B_c_329_n N_A_313_74#_c_890_n 0.0232531f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_356 N_RESET_B_c_330_n N_A_313_74#_c_890_n 0.00245852f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_357 N_RESET_B_c_319_n N_A_313_74#_c_890_n 0.0234271f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_358 N_RESET_B_c_331_n N_A_313_74#_c_891_n 0.00253684f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_359 N_RESET_B_c_332_n N_A_313_74#_c_891_n 0.00819203f $X=5.665 $Y=2.035 $X2=0
+ $Y2=0
cc_360 N_RESET_B_c_333_n N_A_313_74#_c_891_n 0.0158138f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_361 N_RESET_B_c_324_n N_A_313_74#_c_892_n 0.0141476f $X=4.87 $Y=2.24 $X2=0
+ $Y2=0
cc_362 N_RESET_B_c_331_n N_A_313_74#_c_892_n 0.00100516f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_363 N_RESET_B_c_332_n N_A_313_74#_c_892_n 0.00764771f $X=5.665 $Y=2.035 $X2=0
+ $Y2=0
cc_364 N_RESET_B_c_333_n N_A_313_74#_c_892_n 0.00798692f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_365 N_RESET_B_c_336_n N_A_313_74#_c_892_n 0.00688662f $X=5.25 $Y=1.835 $X2=0
+ $Y2=0
cc_366 N_RESET_B_c_331_n N_A_313_74#_c_873_n 0.00690177f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_367 N_RESET_B_c_317_n N_A_699_463#_c_1086_n 0.00129161f $X=4.885 $Y=1.26
+ $X2=0 $Y2=0
cc_368 N_RESET_B_c_331_n N_A_699_463#_c_1095_n 0.00294805f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_369 N_RESET_B_c_332_n N_A_699_463#_c_1095_n 0.00178273f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_370 N_RESET_B_c_333_n N_A_699_463#_c_1095_n 0.00272844f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_371 N_RESET_B_c_315_n N_A_699_463#_c_1087_n 0.00381437f $X=4.885 $Y=1.67
+ $X2=0 $Y2=0
cc_372 N_RESET_B_c_331_n N_A_699_463#_c_1087_n 0.0095029f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_373 N_RESET_B_c_333_n N_A_699_463#_c_1089_n 0.00183407f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_374 N_RESET_B_c_336_n N_A_699_463#_c_1089_n 0.0021429f $X=5.25 $Y=1.835 $X2=0
+ $Y2=0
cc_375 N_RESET_B_c_329_n N_A_699_463#_c_1090_n 0.020213f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_376 N_RESET_B_c_329_n N_A_699_463#_c_1110_n 0.0148124f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_377 N_RESET_B_c_329_n N_A_699_463#_c_1098_n 0.0077093f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_378 N_RESET_B_c_323_n N_A_699_463#_c_1091_n 0.00324495f $X=4.87 $Y=2.15 $X2=0
+ $Y2=0
cc_379 N_RESET_B_c_324_n N_A_699_463#_c_1091_n 0.0064566f $X=4.87 $Y=2.24 $X2=0
+ $Y2=0
cc_380 N_RESET_B_c_315_n N_A_699_463#_c_1091_n 0.0090051f $X=4.885 $Y=1.67 $X2=0
+ $Y2=0
cc_381 N_RESET_B_c_328_n N_A_699_463#_c_1091_n 0.00990343f $X=4.87 $Y=1.835
+ $X2=0 $Y2=0
cc_382 N_RESET_B_c_329_n N_A_699_463#_c_1091_n 0.0210119f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_383 N_RESET_B_c_332_n N_A_699_463#_c_1091_n 0.00123974f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_384 N_RESET_B_c_333_n N_A_699_463#_c_1091_n 0.0325452f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_385 N_RESET_B_c_315_n N_A_699_463#_c_1092_n 0.00273309f $X=4.885 $Y=1.67
+ $X2=0 $Y2=0
cc_386 N_RESET_B_c_317_n N_A_699_463#_c_1092_n 0.0056443f $X=4.885 $Y=1.26 $X2=0
+ $Y2=0
cc_387 N_RESET_B_c_315_n N_A_699_463#_c_1093_n 0.00501004f $X=4.885 $Y=1.67
+ $X2=0 $Y2=0
cc_388 N_RESET_B_c_317_n N_A_699_463#_c_1093_n 0.00303885f $X=4.885 $Y=1.26
+ $X2=0 $Y2=0
cc_389 N_RESET_B_c_329_n N_A_699_463#_c_1093_n 0.0065884f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_390 N_RESET_B_c_331_n N_A_699_463#_c_1093_n 0.0103027f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_391 N_RESET_B_c_332_n N_A_699_463#_c_1093_n 0.0023311f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_392 N_RESET_B_c_333_n N_A_699_463#_c_1093_n 0.0429796f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_393 N_RESET_B_c_336_n N_A_699_463#_c_1093_n 0.0124264f $X=5.25 $Y=1.835 $X2=0
+ $Y2=0
cc_394 N_RESET_B_c_324_n N_A_699_463#_c_1100_n 0.0161824f $X=4.87 $Y=2.24 $X2=0
+ $Y2=0
cc_395 N_RESET_B_c_329_n N_A_699_463#_c_1100_n 0.00889212f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_396 N_RESET_B_c_333_n N_A_699_463#_c_1100_n 0.00739632f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_397 N_RESET_B_c_336_n N_A_699_463#_c_1100_n 0.00440403f $X=5.25 $Y=1.835
+ $X2=0 $Y2=0
cc_398 N_RESET_B_c_326_n N_A_1678_395#_c_1227_n 0.011773f $X=9.02 $Y=2.39 $X2=0
+ $Y2=0
cc_399 N_RESET_B_c_334_n N_A_1678_395#_c_1227_n 3.76177e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_400 N_RESET_B_c_335_n N_A_1678_395#_c_1227_n 0.0011165f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_401 N_RESET_B_c_326_n N_A_1678_395#_c_1228_n 0.0097334f $X=9.02 $Y=2.39 $X2=0
+ $Y2=0
cc_402 N_RESET_B_M1031_g N_A_1678_395#_M1023_g 0.0119923f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_403 N_RESET_B_c_326_n N_A_1678_395#_c_1220_n 0.0114583f $X=9.02 $Y=2.39 $X2=0
+ $Y2=0
cc_404 N_RESET_B_M1031_g N_A_1678_395#_c_1220_n 0.0189876f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_405 N_RESET_B_c_331_n N_A_1678_395#_c_1220_n 0.00170338f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_406 N_RESET_B_c_334_n N_A_1678_395#_c_1220_n 7.09824e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_407 N_RESET_B_c_335_n N_A_1678_395#_c_1220_n 0.00127122f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_408 N_RESET_B_c_331_n N_A_1678_395#_c_1230_n 0.00849993f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_409 N_RESET_B_c_334_n N_A_1678_395#_c_1230_n 3.05552e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_410 N_RESET_B_M1031_g N_A_1678_395#_c_1221_n 0.0151687f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_411 N_RESET_B_c_326_n N_A_1678_395#_c_1231_n 0.00406986f $X=9.02 $Y=2.39
+ $X2=0 $Y2=0
cc_412 N_RESET_B_c_334_n N_A_1678_395#_c_1231_n 5.78327e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_413 N_RESET_B_c_335_n N_A_1678_395#_c_1231_n 0.016871f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_414 N_RESET_B_c_326_n N_A_1678_395#_c_1233_n 3.78573e-19 $X=9.02 $Y=2.39
+ $X2=0 $Y2=0
cc_415 N_RESET_B_M1031_g N_A_1678_395#_c_1233_n 0.00130041f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_416 N_RESET_B_c_334_n N_A_1678_395#_c_1233_n 7.6951e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_417 N_RESET_B_c_335_n N_A_1678_395#_c_1233_n 0.0098343f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_418 N_RESET_B_M1031_g N_A_1678_395#_c_1222_n 0.00227582f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_419 N_RESET_B_M1031_g N_A_1678_395#_c_1224_n 0.00118187f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_420 N_RESET_B_M1031_g N_A_1678_395#_c_1225_n 0.021263f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_421 N_RESET_B_c_326_n N_A_1678_395#_c_1235_n 0.00689999f $X=9.02 $Y=2.39
+ $X2=0 $Y2=0
cc_422 N_RESET_B_c_335_n N_A_1678_395#_c_1235_n 0.00483781f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_423 N_RESET_B_c_331_n N_A_1350_392#_M1011_d 0.00395996f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_424 N_RESET_B_M1031_g N_A_1350_392#_M1032_g 0.0569104f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_425 N_RESET_B_c_326_n N_A_1350_392#_c_1357_n 0.023064f $X=9.02 $Y=2.39 $X2=0
+ $Y2=0
cc_426 N_RESET_B_M1031_g N_A_1350_392#_c_1357_n 0.0128751f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_427 N_RESET_B_c_335_n N_A_1350_392#_c_1357_n 4.39619e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_428 N_RESET_B_c_326_n N_A_1350_392#_c_1358_n 0.00918927f $X=9.02 $Y=2.39
+ $X2=0 $Y2=0
cc_429 N_RESET_B_c_331_n N_A_1350_392#_c_1351_n 0.0218301f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_430 N_RESET_B_c_331_n N_A_1350_392#_c_1380_n 0.0243354f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_431 N_RESET_B_c_326_n N_A_1350_392#_c_1368_n 0.00113733f $X=9.02 $Y=2.39
+ $X2=0 $Y2=0
cc_432 N_RESET_B_c_331_n N_A_1350_392#_c_1368_n 0.023506f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_433 N_RESET_B_c_334_n N_A_1350_392#_c_1368_n 0.00234791f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_434 N_RESET_B_c_335_n N_A_1350_392#_c_1368_n 0.0125499f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_435 N_RESET_B_c_326_n N_A_1350_392#_c_1353_n 0.00113327f $X=9.02 $Y=2.39
+ $X2=0 $Y2=0
cc_436 N_RESET_B_M1031_g N_A_1350_392#_c_1353_n 0.0116508f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_437 N_RESET_B_c_331_n N_A_1350_392#_c_1353_n 0.0123609f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_438 N_RESET_B_c_334_n N_A_1350_392#_c_1353_n 0.00816472f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_439 N_RESET_B_c_335_n N_A_1350_392#_c_1353_n 0.0203289f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_440 N_RESET_B_M1031_g N_A_1350_392#_c_1355_n 0.00118604f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_441 N_RESET_B_M1031_g N_A_1350_392#_c_1356_n 0.0213066f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_442 N_RESET_B_c_329_n N_VPWR_M1004_d 0.00601357f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_443 N_RESET_B_c_331_n N_VPWR_M1005_s 0.00715041f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_444 N_RESET_B_c_322_n N_VPWR_c_1643_n 0.00589882f $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_445 N_RESET_B_c_324_n N_VPWR_c_1645_n 0.00332804f $X=4.87 $Y=2.24 $X2=0 $Y2=0
cc_446 N_RESET_B_c_326_n N_VPWR_c_1647_n 0.00837136f $X=9.02 $Y=2.39 $X2=0 $Y2=0
cc_447 N_RESET_B_c_331_n N_VPWR_c_1647_n 0.00679776f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_448 N_RESET_B_c_334_n N_VPWR_c_1647_n 0.0023649f $X=8.88 $Y=2.035 $X2=0 $Y2=0
cc_449 N_RESET_B_c_335_n N_VPWR_c_1647_n 0.0114656f $X=8.88 $Y=2.035 $X2=0 $Y2=0
cc_450 N_RESET_B_c_326_n N_VPWR_c_1655_n 0.0050971f $X=9.02 $Y=2.39 $X2=0 $Y2=0
cc_451 N_RESET_B_c_322_n N_VPWR_c_1659_n 0.00444469f $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_452 N_RESET_B_c_322_n N_VPWR_c_1640_n 0.0046079f $X=0.95 $Y=2.465 $X2=0 $Y2=0
cc_453 N_RESET_B_c_324_n N_VPWR_c_1640_n 9.39239e-19 $X=4.87 $Y=2.24 $X2=0 $Y2=0
cc_454 N_RESET_B_c_326_n N_VPWR_c_1640_n 0.0052212f $X=9.02 $Y=2.39 $X2=0 $Y2=0
cc_455 N_RESET_B_M1009_g N_A_37_78#_c_1805_n 7.80212e-19 $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_456 N_RESET_B_M1009_g N_A_37_78#_c_1806_n 0.0165609f $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_457 N_RESET_B_c_330_n N_A_37_78#_c_1806_n 0.00197026f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_458 N_RESET_B_c_319_n N_A_37_78#_c_1806_n 0.0729934f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_459 N_RESET_B_c_329_n N_A_37_78#_c_1813_n 0.0300223f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_460 N_RESET_B_c_329_n N_A_37_78#_c_1814_n 0.0173569f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_461 N_RESET_B_c_329_n N_A_37_78#_c_1808_n 0.00328533f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_462 N_RESET_B_c_329_n N_A_37_78#_c_1809_n 5.06485e-19 $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_463 N_RESET_B_c_329_n N_A_37_78#_c_1810_n 0.0103535f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_464 N_RESET_B_M1009_g N_A_37_78#_c_1811_n 8.54775e-19 $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_465 N_RESET_B_c_321_n N_A_37_78#_c_1816_n 0.00220362f $X=0.95 $Y=2.375 $X2=0
+ $Y2=0
cc_466 N_RESET_B_c_322_n N_A_37_78#_c_1816_n 0.012959f $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_467 N_RESET_B_c_321_n N_A_37_78#_c_1817_n 0.00855069f $X=0.95 $Y=2.375 $X2=0
+ $Y2=0
cc_468 N_RESET_B_c_322_n N_A_37_78#_c_1817_n 0.00725597f $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_469 N_RESET_B_c_329_n N_A_37_78#_c_1817_n 0.00640759f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_470 N_RESET_B_c_330_n N_A_37_78#_c_1817_n 0.00929883f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_471 N_RESET_B_c_319_n N_A_37_78#_c_1817_n 0.0168317f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_472 N_RESET_B_c_338_n N_A_37_78#_c_1817_n 0.00290874f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_473 N_RESET_B_c_322_n N_A_37_78#_c_1818_n 5.09312e-19 $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_474 N_RESET_B_c_329_n N_A_37_78#_c_1819_n 0.0212115f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_475 N_RESET_B_M1009_g N_VGND_c_2006_n 0.00582232f $X=0.935 $Y=0.6 $X2=0 $Y2=0
cc_476 N_RESET_B_c_318_n N_VGND_c_2006_n 0.00122895f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_477 N_RESET_B_c_319_n N_VGND_c_2006_n 0.00978084f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_478 N_RESET_B_M1031_g N_VGND_c_2008_n 0.00393134f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_479 N_RESET_B_M1009_g N_VGND_c_2014_n 0.00563421f $X=0.935 $Y=0.6 $X2=0 $Y2=0
cc_480 N_RESET_B_M1031_g N_VGND_c_2016_n 0.00552345f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_481 N_RESET_B_c_314_n N_VGND_c_2019_n 6.39631e-19 $X=4.765 $Y=1.185 $X2=0
+ $Y2=0
cc_482 N_RESET_B_M1009_g N_VGND_c_2029_n 0.00539454f $X=0.935 $Y=0.6 $X2=0 $Y2=0
cc_483 N_RESET_B_M1031_g N_VGND_c_2029_n 0.00534666f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_484 CLK N_A_494_366#_c_576_n 0.003849f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_485 N_CLK_c_527_n N_A_494_366#_c_596_n 0.0013544f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_486 CLK N_A_494_366#_c_596_n 0.00467489f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_487 N_CLK_c_527_n N_A_313_74#_c_874_n 0.0412151f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_488 N_CLK_M1026_g N_A_313_74#_c_859_n 0.0219283f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_489 N_CLK_M1026_g N_A_313_74#_c_865_n 0.00483559f $X=1.925 $Y=0.74 $X2=0
+ $Y2=0
cc_490 N_CLK_c_527_n N_A_313_74#_c_865_n 0.0213194f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_491 CLK N_A_313_74#_c_865_n 0.00554445f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_492 N_CLK_c_527_n N_A_313_74#_c_866_n 0.00475322f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_493 N_CLK_M1026_g N_A_313_74#_c_867_n 0.0101056f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_494 N_CLK_M1026_g N_A_313_74#_c_868_n 0.00364144f $X=1.925 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_CLK_c_527_n N_A_313_74#_c_868_n 0.00484238f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_496 CLK N_A_313_74#_c_868_n 0.031414f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_497 N_CLK_M1026_g N_A_313_74#_c_869_n 0.0117933f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_498 N_CLK_c_527_n N_A_313_74#_c_869_n 6.67273e-19 $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_499 CLK N_A_313_74#_c_869_n 0.0309679f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_500 N_CLK_M1026_g N_A_313_74#_c_870_n 8.37995e-19 $X=1.925 $Y=0.74 $X2=0
+ $Y2=0
cc_501 CLK N_A_313_74#_c_870_n 0.019143f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_502 N_CLK_M1026_g N_A_313_74#_c_872_n 0.00131832f $X=1.925 $Y=0.74 $X2=0
+ $Y2=0
cc_503 N_CLK_c_527_n N_A_313_74#_c_872_n 0.0013406f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_504 CLK N_A_313_74#_c_872_n 0.00666699f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_505 N_CLK_c_527_n N_A_313_74#_c_890_n 0.00404277f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_506 CLK N_A_313_74#_c_890_n 7.47611e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_507 N_CLK_c_527_n N_VPWR_c_1643_n 0.00705047f $X=1.945 $Y=1.755 $X2=0 $Y2=0
cc_508 N_CLK_c_527_n N_VPWR_c_1644_n 0.0106985f $X=1.945 $Y=1.755 $X2=0 $Y2=0
cc_509 N_CLK_c_527_n N_VPWR_c_1660_n 0.00512473f $X=1.945 $Y=1.755 $X2=0 $Y2=0
cc_510 N_CLK_c_527_n N_VPWR_c_1640_n 0.00492022f $X=1.945 $Y=1.755 $X2=0 $Y2=0
cc_511 N_CLK_c_527_n N_A_37_78#_c_1813_n 0.0141735f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_512 CLK N_A_37_78#_c_1813_n 0.00297855f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_513 N_CLK_c_527_n N_A_37_78#_c_1818_n 0.00116669f $X=1.945 $Y=1.755 $X2=0
+ $Y2=0
cc_514 N_CLK_M1026_g N_VGND_c_2006_n 0.00308332f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_515 N_CLK_M1026_g N_VGND_c_2007_n 0.00598308f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_516 N_CLK_M1026_g N_VGND_c_2018_n 0.00434272f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_517 N_CLK_M1026_g N_VGND_c_2029_n 0.00826311f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_518 N_A_494_366#_c_579_n N_A_834_355#_M1017_d 0.0186644f $X=8.105 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_519 N_A_494_366#_c_589_n N_A_834_355#_c_774_n 0.00377028f $X=3.42 $Y=2.15
+ $X2=0 $Y2=0
cc_520 N_A_494_366#_c_588_n N_A_834_355#_c_774_n 0.00121772f $X=3.355 $Y=1.665
+ $X2=0 $Y2=0
cc_521 N_A_494_366#_c_571_n N_A_834_355#_M1025_g 0.00574617f $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_522 N_A_494_366#_M1035_g N_A_834_355#_M1025_g 0.0491928f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_523 N_A_494_366#_c_577_n N_A_834_355#_M1025_g 2.33973e-19 $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_524 N_A_494_366#_c_578_n N_A_834_355#_M1025_g 3.87813e-19 $X=5.395 $Y=0.625
+ $X2=0 $Y2=0
cc_525 N_A_494_366#_c_584_n N_A_834_355#_M1025_g 0.00891123f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_526 N_A_494_366#_M1035_g N_A_834_355#_c_772_n 5.34274e-19 $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_527 N_A_494_366#_c_578_n N_A_834_355#_c_807_n 0.00512559f $X=5.395 $Y=0.625
+ $X2=0 $Y2=0
cc_528 N_A_494_366#_c_584_n N_A_834_355#_c_807_n 0.0116732f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_529 N_A_494_366#_c_579_n N_A_834_355#_c_809_n 0.0530777f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_530 N_A_494_366#_c_578_n N_A_834_355#_c_793_n 0.050878f $X=5.395 $Y=0.625
+ $X2=0 $Y2=0
cc_531 N_A_494_366#_c_579_n N_A_834_355#_c_793_n 0.00379885f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_532 N_A_494_366#_c_585_n N_A_834_355#_c_793_n 0.0123656f $X=5.48 $Y=0.34
+ $X2=0 $Y2=0
cc_533 N_A_494_366#_c_596_n N_A_313_74#_c_874_n 0.00816298f $X=3.015 $Y=1.805
+ $X2=0 $Y2=0
cc_534 N_A_494_366#_c_576_n N_A_313_74#_c_859_n 0.00493406f $X=2.93 $Y=1.72
+ $X2=0 $Y2=0
cc_535 N_A_494_366#_c_582_n N_A_313_74#_c_859_n 0.00714577f $X=2.78 $Y=0.415
+ $X2=0 $Y2=0
cc_536 N_A_494_366#_c_570_n N_A_313_74#_c_860_n 0.00199061f $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_537 N_A_494_366#_c_576_n N_A_313_74#_c_860_n 0.0126774f $X=2.93 $Y=1.72 $X2=0
+ $Y2=0
cc_538 N_A_494_366#_c_595_n N_A_313_74#_c_860_n 0.00472137f $X=3.19 $Y=1.805
+ $X2=0 $Y2=0
cc_539 N_A_494_366#_c_596_n N_A_313_74#_c_860_n 5.85433e-19 $X=3.015 $Y=1.805
+ $X2=0 $Y2=0
cc_540 N_A_494_366#_c_583_n N_A_313_74#_c_860_n 3.05237e-19 $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_541 N_A_494_366#_c_588_n N_A_313_74#_c_860_n 0.0214863f $X=3.355 $Y=1.665
+ $X2=0 $Y2=0
cc_542 N_A_494_366#_c_589_n N_A_313_74#_c_875_n 0.011771f $X=3.42 $Y=2.15 $X2=0
+ $Y2=0
cc_543 N_A_494_366#_c_590_n N_A_313_74#_c_875_n 0.0131071f $X=3.42 $Y=2.24 $X2=0
+ $Y2=0
cc_544 N_A_494_366#_c_596_n N_A_313_74#_c_875_n 0.0172631f $X=3.015 $Y=1.805
+ $X2=0 $Y2=0
cc_545 N_A_494_366#_c_590_n N_A_313_74#_c_876_n 0.0103487f $X=3.42 $Y=2.24 $X2=0
+ $Y2=0
cc_546 N_A_494_366#_M1035_g N_A_313_74#_c_861_n 0.0190138f $X=3.985 $Y=0.9 $X2=0
+ $Y2=0
cc_547 N_A_494_366#_c_577_n N_A_313_74#_c_861_n 0.00661564f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_548 N_A_494_366#_c_582_n N_A_313_74#_c_861_n 0.00459113f $X=2.78 $Y=0.415
+ $X2=0 $Y2=0
cc_549 N_A_494_366#_c_590_n N_A_313_74#_c_878_n 0.00278823f $X=3.42 $Y=2.24
+ $X2=0 $Y2=0
cc_550 N_A_494_366#_c_590_n N_A_313_74#_c_880_n 0.0111333f $X=3.42 $Y=2.24 $X2=0
+ $Y2=0
cc_551 N_A_494_366#_c_570_n N_A_313_74#_c_880_n 0.00457948f $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_494_366#_c_575_n N_A_313_74#_c_862_n 0.00558264f $X=7.185 $Y=1.27
+ $X2=0 $Y2=0
cc_553 N_A_494_366#_c_575_n N_A_313_74#_c_863_n 0.0477631f $X=7.185 $Y=1.27
+ $X2=0 $Y2=0
cc_554 N_A_494_366#_c_593_n N_A_313_74#_c_863_n 0.0233928f $X=8.06 $Y=2.39 $X2=0
+ $Y2=0
cc_555 N_A_494_366#_c_580_n N_A_313_74#_c_863_n 0.0163868f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_556 N_A_494_366#_c_587_n N_A_313_74#_c_863_n 0.0018416f $X=8.19 $Y=1.18 $X2=0
+ $Y2=0
cc_557 N_A_494_366#_c_579_n N_A_313_74#_M1037_g 0.0088085f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_558 N_A_494_366#_c_580_n N_A_313_74#_M1037_g 0.00916962f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_559 N_A_494_366#_c_581_n N_A_313_74#_M1037_g 0.0233298f $X=8.19 $Y=1.015
+ $X2=0 $Y2=0
cc_560 N_A_494_366#_c_586_n N_A_313_74#_M1037_g 0.0213806f $X=7.71 $Y=1.18 $X2=0
+ $Y2=0
cc_561 N_A_494_366#_c_587_n N_A_313_74#_M1037_g 0.0144366f $X=8.19 $Y=1.18 $X2=0
+ $Y2=0
cc_562 N_A_494_366#_c_582_n N_A_313_74#_c_865_n 0.00547313f $X=2.78 $Y=0.415
+ $X2=0 $Y2=0
cc_563 N_A_494_366#_c_576_n N_A_313_74#_c_866_n 0.00526553f $X=2.93 $Y=1.72
+ $X2=0 $Y2=0
cc_564 N_A_494_366#_c_596_n N_A_313_74#_c_866_n 0.0170115f $X=3.015 $Y=1.805
+ $X2=0 $Y2=0
cc_565 N_A_494_366#_c_583_n N_A_313_74#_c_866_n 2.7079e-19 $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_566 N_A_494_366#_c_588_n N_A_313_74#_c_866_n 0.0196386f $X=3.355 $Y=1.665
+ $X2=0 $Y2=0
cc_567 N_A_494_366#_M1012_d N_A_313_74#_c_869_n 0.00207068f $X=2.57 $Y=0.37
+ $X2=0 $Y2=0
cc_568 N_A_494_366#_c_576_n N_A_313_74#_c_869_n 0.0139237f $X=2.93 $Y=1.72 $X2=0
+ $Y2=0
cc_569 N_A_494_366#_c_582_n N_A_313_74#_c_869_n 0.00611482f $X=2.78 $Y=0.415
+ $X2=0 $Y2=0
cc_570 N_A_494_366#_c_576_n N_A_313_74#_c_870_n 0.029587f $X=2.93 $Y=1.72 $X2=0
+ $Y2=0
cc_571 N_A_494_366#_c_596_n N_A_313_74#_c_870_n 0.0169101f $X=3.015 $Y=1.805
+ $X2=0 $Y2=0
cc_572 N_A_494_366#_c_576_n N_A_313_74#_c_871_n 0.00149933f $X=2.93 $Y=1.72
+ $X2=0 $Y2=0
cc_573 N_A_494_366#_c_596_n N_A_313_74#_c_890_n 0.00677034f $X=3.015 $Y=1.805
+ $X2=0 $Y2=0
cc_574 N_A_494_366#_c_575_n N_A_313_74#_c_873_n 7.01297e-19 $X=7.185 $Y=1.27
+ $X2=0 $Y2=0
cc_575 N_A_494_366#_c_579_n N_A_699_463#_c_1086_n 0.013057f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_576 N_A_494_366#_c_585_n N_A_699_463#_c_1086_n 0.00165256f $X=5.48 $Y=0.34
+ $X2=0 $Y2=0
cc_577 N_A_494_366#_c_589_n N_A_699_463#_c_1090_n 4.38636e-19 $X=3.42 $Y=2.15
+ $X2=0 $Y2=0
cc_578 N_A_494_366#_c_571_n N_A_699_463#_c_1090_n 0.00787964f $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_579 N_A_494_366#_M1035_g N_A_699_463#_c_1090_n 0.00704685f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_580 N_A_494_366#_c_590_n N_A_699_463#_c_1098_n 0.00147073f $X=3.42 $Y=2.24
+ $X2=0 $Y2=0
cc_581 N_A_494_366#_c_570_n N_A_699_463#_c_1098_n 0.00117299f $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_582 N_A_494_366#_c_570_n N_A_699_463#_c_1094_n 7.41936e-19 $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_583 N_A_494_366#_c_571_n N_A_699_463#_c_1094_n 0.00282934f $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_584 N_A_494_366#_M1035_g N_A_699_463#_c_1094_n 0.0118197f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_585 N_A_494_366#_c_577_n N_A_699_463#_c_1094_n 0.0325843f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_586 N_A_494_366#_c_584_n N_A_699_463#_c_1094_n 0.00153321f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_587 N_A_494_366#_c_593_n N_A_1678_395#_c_1228_n 0.0291374f $X=8.06 $Y=2.39
+ $X2=0 $Y2=0
cc_588 N_A_494_366#_c_579_n N_A_1678_395#_M1023_g 0.00112332f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_589 N_A_494_366#_c_581_n N_A_1678_395#_M1023_g 0.00454635f $X=8.19 $Y=1.015
+ $X2=0 $Y2=0
cc_590 N_A_494_366#_c_587_n N_A_1678_395#_M1023_g 4.94468e-19 $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_591 N_A_494_366#_c_593_n N_A_1678_395#_c_1230_n 0.0222836f $X=8.06 $Y=2.39
+ $X2=0 $Y2=0
cc_592 N_A_494_366#_c_580_n N_A_1678_395#_c_1230_n 3.41493e-19 $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_593 N_A_494_366#_c_580_n N_A_1678_395#_c_1224_n 8.76782e-19 $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_594 N_A_494_366#_c_587_n N_A_1678_395#_c_1224_n 0.026059f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_595 N_A_494_366#_c_587_n N_A_1678_395#_c_1225_n 0.00189496f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_596 N_A_494_366#_c_579_n N_A_1350_392#_M1006_d 0.00949814f $X=8.105 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_597 N_A_494_366#_c_573_n N_A_1350_392#_c_1393_n 0.00759713f $X=7.11 $Y=1.195
+ $X2=0 $Y2=0
cc_598 N_A_494_366#_c_579_n N_A_1350_392#_c_1393_n 0.00844204f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_599 N_A_494_366#_c_573_n N_A_1350_392#_c_1351_n 0.0120402f $X=7.11 $Y=1.195
+ $X2=0 $Y2=0
cc_600 N_A_494_366#_c_574_n N_A_1350_392#_c_1351_n 0.00910494f $X=7.545 $Y=1.27
+ $X2=0 $Y2=0
cc_601 N_A_494_366#_c_575_n N_A_1350_392#_c_1351_n 0.00382426f $X=7.185 $Y=1.27
+ $X2=0 $Y2=0
cc_602 N_A_494_366#_c_593_n N_A_1350_392#_c_1351_n 0.00895259f $X=8.06 $Y=2.39
+ $X2=0 $Y2=0
cc_603 N_A_494_366#_c_580_n N_A_1350_392#_c_1351_n 0.036911f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_604 N_A_494_366#_c_586_n N_A_1350_392#_c_1351_n 6.23735e-19 $X=7.71 $Y=1.18
+ $X2=0 $Y2=0
cc_605 N_A_494_366#_c_587_n N_A_1350_392#_c_1351_n 0.0212415f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_606 N_A_494_366#_c_574_n N_A_1350_392#_c_1352_n 0.00633476f $X=7.545 $Y=1.27
+ $X2=0 $Y2=0
cc_607 N_A_494_366#_c_579_n N_A_1350_392#_c_1352_n 0.0424696f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_608 N_A_494_366#_c_581_n N_A_1350_392#_c_1352_n 0.0196081f $X=8.19 $Y=1.015
+ $X2=0 $Y2=0
cc_609 N_A_494_366#_c_586_n N_A_1350_392#_c_1352_n 0.00746605f $X=7.71 $Y=1.18
+ $X2=0 $Y2=0
cc_610 N_A_494_366#_c_587_n N_A_1350_392#_c_1352_n 0.030444f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_611 N_A_494_366#_c_593_n N_A_1350_392#_c_1380_n 0.014773f $X=8.06 $Y=2.39
+ $X2=0 $Y2=0
cc_612 N_A_494_366#_c_580_n N_A_1350_392#_c_1380_n 0.0233132f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_613 N_A_494_366#_c_593_n N_A_1350_392#_c_1368_n 0.00585809f $X=8.06 $Y=2.39
+ $X2=0 $Y2=0
cc_614 N_A_494_366#_c_580_n N_A_1350_392#_c_1368_n 0.045021f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_615 N_A_494_366#_c_580_n N_A_1350_392#_c_1354_n 0.0145381f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_616 N_A_494_366#_c_587_n N_A_1350_392#_c_1354_n 0.00286183f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_617 N_A_494_366#_c_593_n N_VPWR_c_1653_n 0.00391396f $X=8.06 $Y=2.39 $X2=0
+ $Y2=0
cc_618 N_A_494_366#_c_590_n N_VPWR_c_1640_n 9.39239e-19 $X=3.42 $Y=2.24 $X2=0
+ $Y2=0
cc_619 N_A_494_366#_c_593_n N_VPWR_c_1640_n 0.0052212f $X=8.06 $Y=2.39 $X2=0
+ $Y2=0
cc_620 N_A_494_366#_M1010_d N_A_37_78#_c_1813_n 0.00655641f $X=2.47 $Y=1.83
+ $X2=0 $Y2=0
cc_621 N_A_494_366#_c_595_n N_A_37_78#_c_1813_n 2.61867e-19 $X=3.19 $Y=1.805
+ $X2=0 $Y2=0
cc_622 N_A_494_366#_c_596_n N_A_37_78#_c_1813_n 0.0271291f $X=3.015 $Y=1.805
+ $X2=0 $Y2=0
cc_623 N_A_494_366#_M1035_g N_A_37_78#_c_1807_n 6.83611e-19 $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_624 N_A_494_366#_c_577_n N_A_37_78#_c_1807_n 0.0198813f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_625 N_A_494_366#_c_582_n N_A_37_78#_c_1807_n 0.043075f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_626 N_A_494_366#_c_589_n N_A_37_78#_c_1814_n 0.00457619f $X=3.42 $Y=2.15
+ $X2=0 $Y2=0
cc_627 N_A_494_366#_c_590_n N_A_37_78#_c_1814_n 0.00875594f $X=3.42 $Y=2.24
+ $X2=0 $Y2=0
cc_628 N_A_494_366#_c_570_n N_A_37_78#_c_1814_n 0.00189986f $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_629 N_A_494_366#_c_583_n N_A_37_78#_c_1814_n 0.00585052f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_630 N_A_494_366#_c_588_n N_A_37_78#_c_1814_n 2.58281e-19 $X=3.355 $Y=1.665
+ $X2=0 $Y2=0
cc_631 N_A_494_366#_c_570_n N_A_37_78#_c_1808_n 0.0018714f $X=3.8 $Y=1.665 $X2=0
+ $Y2=0
cc_632 N_A_494_366#_M1035_g N_A_37_78#_c_1808_n 0.00174133f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_633 N_A_494_366#_c_583_n N_A_37_78#_c_1808_n 0.00136135f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_634 N_A_494_366#_c_588_n N_A_37_78#_c_1808_n 7.58999e-19 $X=3.355 $Y=1.665
+ $X2=0 $Y2=0
cc_635 N_A_494_366#_c_576_n N_A_37_78#_c_1809_n 0.0131612f $X=2.93 $Y=1.72 $X2=0
+ $Y2=0
cc_636 N_A_494_366#_c_595_n N_A_37_78#_c_1809_n 2.34784e-19 $X=3.19 $Y=1.805
+ $X2=0 $Y2=0
cc_637 N_A_494_366#_c_583_n N_A_37_78#_c_1809_n 0.0201764f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_638 N_A_494_366#_c_588_n N_A_37_78#_c_1809_n 9.19535e-19 $X=3.355 $Y=1.665
+ $X2=0 $Y2=0
cc_639 N_A_494_366#_c_589_n N_A_37_78#_c_1810_n 0.00398592f $X=3.42 $Y=2.15
+ $X2=0 $Y2=0
cc_640 N_A_494_366#_c_570_n N_A_37_78#_c_1810_n 0.0129932f $X=3.8 $Y=1.665 $X2=0
+ $Y2=0
cc_641 N_A_494_366#_c_571_n N_A_37_78#_c_1810_n 0.00458963f $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_642 N_A_494_366#_c_576_n N_A_37_78#_c_1810_n 0.00524765f $X=2.93 $Y=1.72
+ $X2=0 $Y2=0
cc_643 N_A_494_366#_c_583_n N_A_37_78#_c_1810_n 0.0238297f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_644 N_A_494_366#_c_588_n N_A_37_78#_c_1810_n 0.00239679f $X=3.355 $Y=1.665
+ $X2=0 $Y2=0
cc_645 N_A_494_366#_c_589_n N_A_37_78#_c_1819_n 0.00165814f $X=3.42 $Y=2.15
+ $X2=0 $Y2=0
cc_646 N_A_494_366#_c_590_n N_A_37_78#_c_1819_n 0.0102679f $X=3.42 $Y=2.24 $X2=0
+ $Y2=0
cc_647 N_A_494_366#_c_595_n N_A_37_78#_c_1819_n 0.0106104f $X=3.19 $Y=1.805
+ $X2=0 $Y2=0
cc_648 N_A_494_366#_c_596_n N_A_37_78#_c_1819_n 0.00775205f $X=3.015 $Y=1.805
+ $X2=0 $Y2=0
cc_649 N_A_494_366#_c_583_n N_A_37_78#_c_1819_n 0.0111562f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_650 N_A_494_366#_c_588_n N_A_37_78#_c_1819_n 9.62291e-19 $X=3.355 $Y=1.665
+ $X2=0 $Y2=0
cc_651 N_A_494_366#_c_578_n N_VGND_M1034_d 0.0148411f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_652 N_A_494_366#_c_585_n N_VGND_M1034_d 0.0100088f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_653 N_A_494_366#_c_582_n N_VGND_c_2007_n 0.0202383f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_654 N_A_494_366#_c_579_n N_VGND_c_2008_n 0.00808546f $X=8.105 $Y=0.34 $X2=0
+ $Y2=0
cc_655 N_A_494_366#_c_581_n N_VGND_c_2008_n 0.0105982f $X=8.19 $Y=1.015 $X2=0
+ $Y2=0
cc_656 N_A_494_366#_c_577_n N_VGND_c_2019_n 0.0565209f $X=4.305 $Y=0.415 $X2=0
+ $Y2=0
cc_657 N_A_494_366#_c_578_n N_VGND_c_2019_n 0.00950268f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_658 N_A_494_366#_c_582_n N_VGND_c_2019_n 0.0222466f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_659 N_A_494_366#_c_584_n N_VGND_c_2019_n 0.00781472f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_660 N_A_494_366#_c_573_n N_VGND_c_2020_n 0.00278271f $X=7.11 $Y=1.195 $X2=0
+ $Y2=0
cc_661 N_A_494_366#_c_578_n N_VGND_c_2020_n 0.00371184f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_662 N_A_494_366#_c_579_n N_VGND_c_2020_n 0.174907f $X=8.105 $Y=0.34 $X2=0
+ $Y2=0
cc_663 N_A_494_366#_c_585_n N_VGND_c_2020_n 0.0116868f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_664 N_A_494_366#_c_578_n N_VGND_c_2025_n 0.0242401f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_665 N_A_494_366#_c_584_n N_VGND_c_2025_n 0.00169795f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_666 N_A_494_366#_c_585_n N_VGND_c_2025_n 0.00911753f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_667 N_A_494_366#_c_573_n N_VGND_c_2029_n 0.00363426f $X=7.11 $Y=1.195 $X2=0
+ $Y2=0
cc_668 N_A_494_366#_c_577_n N_VGND_c_2029_n 0.0462418f $X=4.305 $Y=0.415 $X2=0
+ $Y2=0
cc_669 N_A_494_366#_c_578_n N_VGND_c_2029_n 0.0200036f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_670 N_A_494_366#_c_579_n N_VGND_c_2029_n 0.100739f $X=8.105 $Y=0.34 $X2=0
+ $Y2=0
cc_671 N_A_494_366#_c_582_n N_VGND_c_2029_n 0.0172447f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_672 N_A_494_366#_c_584_n N_VGND_c_2029_n 0.00616507f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_673 N_A_494_366#_c_585_n N_VGND_c_2029_n 0.00646475f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_674 N_A_494_366#_c_578_n A_890_138# 0.00133041f $X=5.395 $Y=0.625 $X2=-0.19
+ $Y2=-0.245
cc_675 N_A_834_355#_c_774_n N_A_313_74#_c_878_n 0.0032308f $X=4.26 $Y=2.24 $X2=0
+ $Y2=0
cc_676 N_A_834_355#_c_774_n N_A_313_74#_c_880_n 0.0320057f $X=4.26 $Y=2.24 $X2=0
+ $Y2=0
cc_677 N_A_834_355#_c_774_n N_A_313_74#_c_881_n 0.00995786f $X=4.26 $Y=2.24
+ $X2=0 $Y2=0
cc_678 N_A_834_355#_c_773_n N_A_313_74#_c_862_n 0.0037176f $X=6.24 $Y=1.94 $X2=0
+ $Y2=0
cc_679 N_A_834_355#_c_817_p N_A_313_74#_c_862_n 0.00809783f $X=6.825 $Y=0.885
+ $X2=0 $Y2=0
cc_680 N_A_834_355#_c_778_n N_A_313_74#_c_862_n 0.00544466f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_681 N_A_834_355#_c_817_p N_A_313_74#_c_863_n 8.72478e-19 $X=6.825 $Y=0.885
+ $X2=0 $Y2=0
cc_682 N_A_834_355#_M1005_d N_A_313_74#_c_888_n 0.00553679f $X=6.3 $Y=1.96 $X2=0
+ $Y2=0
cc_683 N_A_834_355#_c_778_n N_A_313_74#_c_888_n 0.0236327f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_684 N_A_834_355#_c_773_n N_A_313_74#_c_889_n 0.0126354f $X=6.24 $Y=1.94 $X2=0
+ $Y2=0
cc_685 N_A_834_355#_c_778_n N_A_313_74#_c_889_n 0.0138472f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_686 N_A_834_355#_c_773_n N_A_313_74#_c_873_n 0.0254145f $X=6.24 $Y=1.94 $X2=0
+ $Y2=0
cc_687 N_A_834_355#_c_817_p N_A_313_74#_c_873_n 0.0309014f $X=6.825 $Y=0.885
+ $X2=0 $Y2=0
cc_688 N_A_834_355#_c_778_n N_A_313_74#_c_873_n 0.00458428f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_689 N_A_834_355#_c_773_n N_A_699_463#_c_1086_n 0.00417334f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_690 N_A_834_355#_c_809_n N_A_699_463#_c_1086_n 0.00865527f $X=6.325 $Y=0.885
+ $X2=0 $Y2=0
cc_691 N_A_834_355#_c_793_n N_A_699_463#_c_1086_n 0.010622f $X=5.735 $Y=0.885
+ $X2=0 $Y2=0
cc_692 N_A_834_355#_c_773_n N_A_699_463#_c_1095_n 0.00803887f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_693 N_A_834_355#_c_778_n N_A_699_463#_c_1095_n 0.011835f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_694 N_A_834_355#_c_773_n N_A_699_463#_c_1088_n 0.0135266f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_695 N_A_834_355#_c_809_n N_A_699_463#_c_1088_n 0.0125467f $X=6.325 $Y=0.885
+ $X2=0 $Y2=0
cc_696 N_A_834_355#_c_773_n N_A_699_463#_c_1089_n 0.00813214f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_697 N_A_834_355#_c_774_n N_A_699_463#_c_1090_n 0.00749506f $X=4.26 $Y=2.24
+ $X2=0 $Y2=0
cc_698 N_A_834_355#_M1025_g N_A_699_463#_c_1090_n 0.00448986f $X=4.375 $Y=0.9
+ $X2=0 $Y2=0
cc_699 N_A_834_355#_c_772_n N_A_699_463#_c_1090_n 0.0773505f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_700 N_A_834_355#_c_774_n N_A_699_463#_c_1110_n 0.0137776f $X=4.26 $Y=2.24
+ $X2=0 $Y2=0
cc_701 N_A_834_355#_c_772_n N_A_699_463#_c_1110_n 0.00796644f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_702 N_A_834_355#_c_774_n N_A_699_463#_c_1098_n 8.75103e-19 $X=4.26 $Y=2.24
+ $X2=0 $Y2=0
cc_703 N_A_834_355#_c_774_n N_A_699_463#_c_1091_n 0.00306279f $X=4.26 $Y=2.24
+ $X2=0 $Y2=0
cc_704 N_A_834_355#_M1025_g N_A_699_463#_c_1091_n 6.92887e-19 $X=4.375 $Y=0.9
+ $X2=0 $Y2=0
cc_705 N_A_834_355#_c_772_n N_A_699_463#_c_1091_n 0.0439058f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_706 N_A_834_355#_M1025_g N_A_699_463#_c_1092_n 6.42461e-19 $X=4.375 $Y=0.9
+ $X2=0 $Y2=0
cc_707 N_A_834_355#_c_772_n N_A_699_463#_c_1092_n 0.0233608f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_708 N_A_834_355#_c_793_n N_A_699_463#_c_1092_n 0.0110525f $X=5.735 $Y=0.885
+ $X2=0 $Y2=0
cc_709 N_A_834_355#_c_773_n N_A_699_463#_c_1093_n 0.0211767f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_710 N_A_834_355#_c_793_n N_A_699_463#_c_1093_n 0.0767028f $X=5.735 $Y=0.885
+ $X2=0 $Y2=0
cc_711 N_A_834_355#_M1025_g N_A_699_463#_c_1094_n 0.00193581f $X=4.375 $Y=0.9
+ $X2=0 $Y2=0
cc_712 N_A_834_355#_c_807_n N_A_699_463#_c_1094_n 0.0145807f $X=4.57 $Y=0.965
+ $X2=0 $Y2=0
cc_713 N_A_834_355#_c_774_n N_A_699_463#_c_1100_n 0.00122425f $X=4.26 $Y=2.24
+ $X2=0 $Y2=0
cc_714 N_A_834_355#_c_774_n N_VPWR_c_1645_n 0.00341428f $X=4.26 $Y=2.24 $X2=0
+ $Y2=0
cc_715 N_A_834_355#_c_774_n N_VPWR_c_1640_n 9.39239e-19 $X=4.26 $Y=2.24 $X2=0
+ $Y2=0
cc_716 N_A_834_355#_c_793_n N_VGND_M1034_d 0.017178f $X=5.735 $Y=0.885 $X2=0
+ $Y2=0
cc_717 N_A_834_355#_M1025_g N_VGND_c_2019_n 5.26406e-19 $X=4.375 $Y=0.9 $X2=0
+ $Y2=0
cc_718 N_A_834_355#_c_772_n A_890_138# 7.01113e-19 $X=4.405 $Y=1.94 $X2=-0.19
+ $Y2=-0.245
cc_719 N_A_834_355#_c_807_n A_890_138# 6.98889e-19 $X=4.57 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_720 N_A_834_355#_c_793_n A_890_138# 0.00302632f $X=5.735 $Y=0.885 $X2=-0.19
+ $Y2=-0.245
cc_721 N_A_313_74#_c_882_n N_A_699_463#_c_1095_n 0.00530352f $X=5.385 $Y=3.075
+ $X2=0 $Y2=0
cc_722 N_A_313_74#_c_862_n N_A_699_463#_c_1095_n 0.0432171f $X=6.675 $Y=1.885
+ $X2=0 $Y2=0
cc_723 N_A_313_74#_c_888_n N_A_699_463#_c_1095_n 0.012815f $X=6.785 $Y=2.49
+ $X2=0 $Y2=0
cc_724 N_A_313_74#_c_891_n N_A_699_463#_c_1095_n 7.70919e-19 $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_725 N_A_313_74#_c_892_n N_A_699_463#_c_1095_n 0.00992481f $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_726 N_A_313_74#_c_892_n N_A_699_463#_c_1087_n 0.00125125f $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_727 N_A_313_74#_c_862_n N_A_699_463#_c_1088_n 0.0214503f $X=6.675 $Y=1.885
+ $X2=0 $Y2=0
cc_728 N_A_313_74#_c_873_n N_A_699_463#_c_1088_n 3.74234e-19 $X=6.87 $Y=1.425
+ $X2=0 $Y2=0
cc_729 N_A_313_74#_c_862_n N_A_699_463#_c_1089_n 0.00590001f $X=6.675 $Y=1.885
+ $X2=0 $Y2=0
cc_730 N_A_313_74#_c_861_n N_A_699_463#_c_1090_n 4.36892e-19 $X=3.485 $Y=1.2
+ $X2=0 $Y2=0
cc_731 N_A_313_74#_c_880_n N_A_699_463#_c_1090_n 0.00150894f $X=3.87 $Y=2.81
+ $X2=0 $Y2=0
cc_732 N_A_313_74#_c_881_n N_A_699_463#_c_1110_n 0.0025284f $X=5.31 $Y=3.15
+ $X2=0 $Y2=0
cc_733 N_A_313_74#_c_876_n N_A_699_463#_c_1098_n 0.00252649f $X=3.78 $Y=3.15
+ $X2=0 $Y2=0
cc_734 N_A_313_74#_c_878_n N_A_699_463#_c_1098_n 4.86419e-19 $X=3.87 $Y=2.9
+ $X2=0 $Y2=0
cc_735 N_A_313_74#_c_880_n N_A_699_463#_c_1098_n 0.0123709f $X=3.87 $Y=2.81
+ $X2=0 $Y2=0
cc_736 N_A_313_74#_c_881_n N_A_699_463#_c_1098_n 0.00145066f $X=5.31 $Y=3.15
+ $X2=0 $Y2=0
cc_737 N_A_313_74#_c_892_n N_A_699_463#_c_1091_n 5.20942e-19 $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_738 N_A_313_74#_c_861_n N_A_699_463#_c_1094_n 0.00204771f $X=3.485 $Y=1.2
+ $X2=0 $Y2=0
cc_739 N_A_313_74#_c_881_n N_A_699_463#_c_1100_n 0.00497916f $X=5.31 $Y=3.15
+ $X2=0 $Y2=0
cc_740 N_A_313_74#_c_891_n N_A_699_463#_c_1100_n 0.0190155f $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_741 N_A_313_74#_c_892_n N_A_699_463#_c_1100_n 0.00698712f $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_742 N_A_313_74#_M1037_g N_A_1678_395#_M1023_g 0.0378955f $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_743 N_A_313_74#_c_863_n N_A_1678_395#_c_1220_n 0.0216911f $X=8.085 $Y=1.66
+ $X2=0 $Y2=0
cc_744 N_A_313_74#_M1037_g N_A_1678_395#_c_1224_n 4.34985e-19 $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_745 N_A_313_74#_M1037_g N_A_1678_395#_c_1225_n 0.0216911f $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_746 N_A_313_74#_c_888_n N_A_1350_392#_M1011_d 0.00523037f $X=6.785 $Y=2.49
+ $X2=0 $Y2=0
cc_747 N_A_313_74#_c_889_n N_A_1350_392#_M1011_d 0.00670815f $X=6.87 $Y=2.405
+ $X2=0 $Y2=0
cc_748 N_A_313_74#_c_862_n N_A_1350_392#_c_1351_n 0.0104964f $X=6.675 $Y=1.885
+ $X2=0 $Y2=0
cc_749 N_A_313_74#_c_863_n N_A_1350_392#_c_1351_n 0.013648f $X=8.085 $Y=1.66
+ $X2=0 $Y2=0
cc_750 N_A_313_74#_c_888_n N_A_1350_392#_c_1351_n 0.0140223f $X=6.785 $Y=2.49
+ $X2=0 $Y2=0
cc_751 N_A_313_74#_c_889_n N_A_1350_392#_c_1351_n 0.0510782f $X=6.87 $Y=2.405
+ $X2=0 $Y2=0
cc_752 N_A_313_74#_c_873_n N_A_1350_392#_c_1351_n 0.0231503f $X=6.87 $Y=1.425
+ $X2=0 $Y2=0
cc_753 N_A_313_74#_M1037_g N_A_1350_392#_c_1352_n 0.00507341f $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_754 N_A_313_74#_c_863_n N_A_1350_392#_c_1368_n 2.44969e-19 $X=8.085 $Y=1.66
+ $X2=0 $Y2=0
cc_755 N_A_313_74#_M1037_g N_A_1350_392#_c_1354_n 0.00153073f $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_756 N_A_313_74#_c_888_n N_VPWR_M1005_s 0.00587787f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_757 N_A_313_74#_c_874_n N_VPWR_c_1644_n 0.0095685f $X=2.395 $Y=1.755 $X2=0
+ $Y2=0
cc_758 N_A_313_74#_c_875_n N_VPWR_c_1644_n 0.00185176f $X=2.905 $Y=3.075 $X2=0
+ $Y2=0
cc_759 N_A_313_74#_c_877_n N_VPWR_c_1644_n 0.00261603f $X=2.98 $Y=3.15 $X2=0
+ $Y2=0
cc_760 N_A_313_74#_c_878_n N_VPWR_c_1645_n 0.00604173f $X=3.87 $Y=2.9 $X2=0
+ $Y2=0
cc_761 N_A_313_74#_c_881_n N_VPWR_c_1645_n 0.0250293f $X=5.31 $Y=3.15 $X2=0
+ $Y2=0
cc_762 N_A_313_74#_c_882_n N_VPWR_c_1645_n 0.00529928f $X=5.385 $Y=3.075 $X2=0
+ $Y2=0
cc_763 N_A_313_74#_c_882_n N_VPWR_c_1646_n 0.0102081f $X=5.385 $Y=3.075 $X2=0
+ $Y2=0
cc_764 N_A_313_74#_c_862_n N_VPWR_c_1646_n 0.00165063f $X=6.675 $Y=1.885 $X2=0
+ $Y2=0
cc_765 N_A_313_74#_c_888_n N_VPWR_c_1646_n 0.0217061f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_766 N_A_313_74#_c_862_n N_VPWR_c_1653_n 0.00338554f $X=6.675 $Y=1.885 $X2=0
+ $Y2=0
cc_767 N_A_313_74#_c_888_n N_VPWR_c_1653_n 0.00955729f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_768 N_A_313_74#_c_874_n N_VPWR_c_1661_n 0.00512473f $X=2.395 $Y=1.755 $X2=0
+ $Y2=0
cc_769 N_A_313_74#_c_877_n N_VPWR_c_1661_n 0.0453861f $X=2.98 $Y=3.15 $X2=0
+ $Y2=0
cc_770 N_A_313_74#_c_881_n N_VPWR_c_1662_n 0.0212613f $X=5.31 $Y=3.15 $X2=0
+ $Y2=0
cc_771 N_A_313_74#_c_888_n N_VPWR_c_1662_n 0.00150121f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_772 N_A_313_74#_c_891_n N_VPWR_c_1662_n 0.00478946f $X=5.56 $Y=2.375 $X2=0
+ $Y2=0
cc_773 N_A_313_74#_c_874_n N_VPWR_c_1640_n 0.00492022f $X=2.395 $Y=1.755 $X2=0
+ $Y2=0
cc_774 N_A_313_74#_c_876_n N_VPWR_c_1640_n 0.0239748f $X=3.78 $Y=3.15 $X2=0
+ $Y2=0
cc_775 N_A_313_74#_c_877_n N_VPWR_c_1640_n 0.00710688f $X=2.98 $Y=3.15 $X2=0
+ $Y2=0
cc_776 N_A_313_74#_c_881_n N_VPWR_c_1640_n 0.0415621f $X=5.31 $Y=3.15 $X2=0
+ $Y2=0
cc_777 N_A_313_74#_c_862_n N_VPWR_c_1640_n 0.00448618f $X=6.675 $Y=1.885 $X2=0
+ $Y2=0
cc_778 N_A_313_74#_c_886_n N_VPWR_c_1640_n 0.00539862f $X=3.87 $Y=3.15 $X2=0
+ $Y2=0
cc_779 N_A_313_74#_c_888_n N_VPWR_c_1640_n 0.0234322f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_780 N_A_313_74#_c_891_n N_VPWR_c_1640_n 0.00841698f $X=5.56 $Y=2.375 $X2=0
+ $Y2=0
cc_781 N_A_313_74#_c_867_n N_A_37_78#_c_1806_n 0.00463142f $X=1.71 $Y=0.515
+ $X2=0 $Y2=0
cc_782 N_A_313_74#_c_872_n N_A_37_78#_c_1806_n 0.00555565f $X=1.665 $Y=1.055
+ $X2=0 $Y2=0
cc_783 N_A_313_74#_M1004_s N_A_37_78#_c_1813_n 0.00410671f $X=1.58 $Y=1.83 $X2=0
+ $Y2=0
cc_784 N_A_313_74#_c_874_n N_A_37_78#_c_1813_n 0.0125528f $X=2.395 $Y=1.755
+ $X2=0 $Y2=0
cc_785 N_A_313_74#_c_875_n N_A_37_78#_c_1813_n 0.0125853f $X=2.905 $Y=3.075
+ $X2=0 $Y2=0
cc_786 N_A_313_74#_c_866_n N_A_37_78#_c_1813_n 9.6488e-19 $X=2.515 $Y=1.59 $X2=0
+ $Y2=0
cc_787 N_A_313_74#_c_890_n N_A_37_78#_c_1813_n 0.00758195f $X=1.72 $Y=1.975
+ $X2=0 $Y2=0
cc_788 N_A_313_74#_c_859_n N_A_37_78#_c_1807_n 9.12798e-19 $X=2.495 $Y=1.2 $X2=0
+ $Y2=0
cc_789 N_A_313_74#_c_860_n N_A_37_78#_c_1807_n 0.0040547f $X=3.41 $Y=1.275 $X2=0
+ $Y2=0
cc_790 N_A_313_74#_c_861_n N_A_37_78#_c_1807_n 0.00939525f $X=3.485 $Y=1.2 $X2=0
+ $Y2=0
cc_791 N_A_313_74#_c_880_n N_A_37_78#_c_1814_n 3.91161e-19 $X=3.87 $Y=2.81 $X2=0
+ $Y2=0
cc_792 N_A_313_74#_c_860_n N_A_37_78#_c_1808_n 0.00854611f $X=3.41 $Y=1.275
+ $X2=0 $Y2=0
cc_793 N_A_313_74#_c_860_n N_A_37_78#_c_1809_n 0.00560277f $X=3.41 $Y=1.275
+ $X2=0 $Y2=0
cc_794 N_A_313_74#_c_890_n N_A_37_78#_c_1817_n 0.016143f $X=1.72 $Y=1.975 $X2=0
+ $Y2=0
cc_795 N_A_313_74#_M1004_s N_A_37_78#_c_1818_n 0.00449636f $X=1.58 $Y=1.83 $X2=0
+ $Y2=0
cc_796 N_A_313_74#_c_875_n N_A_37_78#_c_1819_n 0.0131474f $X=2.905 $Y=3.075
+ $X2=0 $Y2=0
cc_797 N_A_313_74#_c_876_n N_A_37_78#_c_1819_n 0.00561301f $X=3.78 $Y=3.15 $X2=0
+ $Y2=0
cc_798 N_A_313_74#_c_880_n N_A_37_78#_c_1819_n 6.87403e-19 $X=3.87 $Y=2.81 $X2=0
+ $Y2=0
cc_799 N_A_313_74#_c_869_n N_VGND_M1026_d 0.00371446f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_800 N_A_313_74#_c_867_n N_VGND_c_2006_n 0.0317976f $X=1.71 $Y=0.515 $X2=0
+ $Y2=0
cc_801 N_A_313_74#_c_859_n N_VGND_c_2007_n 0.00558618f $X=2.495 $Y=1.2 $X2=0
+ $Y2=0
cc_802 N_A_313_74#_c_867_n N_VGND_c_2007_n 0.0183102f $X=1.71 $Y=0.515 $X2=0
+ $Y2=0
cc_803 N_A_313_74#_c_869_n N_VGND_c_2007_n 0.0248957f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_804 N_A_313_74#_c_867_n N_VGND_c_2018_n 0.0185798f $X=1.71 $Y=0.515 $X2=0
+ $Y2=0
cc_805 N_A_313_74#_c_859_n N_VGND_c_2019_n 0.00433834f $X=2.495 $Y=1.2 $X2=0
+ $Y2=0
cc_806 N_A_313_74#_M1037_g N_VGND_c_2020_n 9.33926e-19 $X=8.16 $Y=0.615 $X2=0
+ $Y2=0
cc_807 N_A_313_74#_c_859_n N_VGND_c_2029_n 0.00826005f $X=2.495 $Y=1.2 $X2=0
+ $Y2=0
cc_808 N_A_313_74#_c_867_n N_VGND_c_2029_n 0.0153224f $X=1.71 $Y=0.515 $X2=0
+ $Y2=0
cc_809 N_A_699_463#_c_1110_n N_VPWR_M1019_d 0.00851579f $X=4.745 $Y=2.485 $X2=0
+ $Y2=0
cc_810 N_A_699_463#_c_1110_n N_VPWR_c_1645_n 0.025965f $X=4.745 $Y=2.485 $X2=0
+ $Y2=0
cc_811 N_A_699_463#_c_1098_n N_VPWR_c_1645_n 4.52709e-19 $X=4.135 $Y=2.485 $X2=0
+ $Y2=0
cc_812 N_A_699_463#_c_1100_n N_VPWR_c_1645_n 0.00110156f $X=4.83 $Y=2.525 $X2=0
+ $Y2=0
cc_813 N_A_699_463#_c_1095_n N_VPWR_c_1646_n 0.00879102f $X=6.225 $Y=1.885 $X2=0
+ $Y2=0
cc_814 N_A_699_463#_c_1100_n N_VPWR_c_1646_n 3.02124e-19 $X=4.83 $Y=2.525 $X2=0
+ $Y2=0
cc_815 N_A_699_463#_c_1095_n N_VPWR_c_1653_n 0.00304117f $X=6.225 $Y=1.885 $X2=0
+ $Y2=0
cc_816 N_A_699_463#_c_1110_n N_VPWR_c_1661_n 0.0027208f $X=4.745 $Y=2.485 $X2=0
+ $Y2=0
cc_817 N_A_699_463#_c_1098_n N_VPWR_c_1661_n 0.00947916f $X=4.135 $Y=2.485 $X2=0
+ $Y2=0
cc_818 N_A_699_463#_c_1100_n N_VPWR_c_1662_n 0.00785197f $X=4.83 $Y=2.525 $X2=0
+ $Y2=0
cc_819 N_A_699_463#_c_1095_n N_VPWR_c_1640_n 0.00395322f $X=6.225 $Y=1.885 $X2=0
+ $Y2=0
cc_820 N_A_699_463#_c_1110_n N_VPWR_c_1640_n 0.00725677f $X=4.745 $Y=2.485 $X2=0
+ $Y2=0
cc_821 N_A_699_463#_c_1098_n N_VPWR_c_1640_n 0.0139664f $X=4.135 $Y=2.485 $X2=0
+ $Y2=0
cc_822 N_A_699_463#_c_1100_n N_VPWR_c_1640_n 0.0110612f $X=4.83 $Y=2.525 $X2=0
+ $Y2=0
cc_823 N_A_699_463#_c_1090_n N_A_37_78#_c_1807_n 0.00327469f $X=4.05 $Y=2.4
+ $X2=0 $Y2=0
cc_824 N_A_699_463#_c_1094_n N_A_37_78#_c_1807_n 0.014524f $X=3.77 $Y=0.86 $X2=0
+ $Y2=0
cc_825 N_A_699_463#_c_1090_n N_A_37_78#_c_1814_n 0.0132299f $X=4.05 $Y=2.4 $X2=0
+ $Y2=0
cc_826 N_A_699_463#_c_1098_n N_A_37_78#_c_1814_n 0.0166624f $X=4.135 $Y=2.485
+ $X2=0 $Y2=0
cc_827 N_A_699_463#_c_1090_n N_A_37_78#_c_1808_n 0.0135526f $X=4.05 $Y=2.4 $X2=0
+ $Y2=0
cc_828 N_A_699_463#_c_1094_n N_A_37_78#_c_1808_n 0.0160421f $X=3.77 $Y=0.86
+ $X2=0 $Y2=0
cc_829 N_A_699_463#_c_1090_n N_A_37_78#_c_1810_n 0.0488054f $X=4.05 $Y=2.4 $X2=0
+ $Y2=0
cc_830 N_A_699_463#_c_1090_n N_A_37_78#_c_1819_n 0.00286442f $X=4.05 $Y=2.4
+ $X2=0 $Y2=0
cc_831 N_A_699_463#_c_1098_n N_A_37_78#_c_1819_n 0.0248711f $X=4.135 $Y=2.485
+ $X2=0 $Y2=0
cc_832 N_A_699_463#_c_1098_n A_789_463# 0.00233332f $X=4.135 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_833 N_A_699_463#_c_1086_n N_VGND_c_2020_n 0.00278271f $X=5.685 $Y=1.22 $X2=0
+ $Y2=0
cc_834 N_A_699_463#_c_1086_n N_VGND_c_2025_n 4.07279e-19 $X=5.685 $Y=1.22 $X2=0
+ $Y2=0
cc_835 N_A_699_463#_c_1086_n N_VGND_c_2029_n 0.00363426f $X=5.685 $Y=1.22 $X2=0
+ $Y2=0
cc_836 N_A_699_463#_c_1090_n A_812_138# 5.10806e-19 $X=4.05 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_837 N_A_699_463#_c_1094_n A_812_138# 0.00174073f $X=3.77 $Y=0.86 $X2=-0.19
+ $Y2=-0.245
cc_838 N_A_1678_395#_c_1221_n N_A_1350_392#_M1032_g 0.0108485f $X=9.5 $Y=1.12
+ $X2=0 $Y2=0
cc_839 N_A_1678_395#_c_1222_n N_A_1350_392#_M1032_g 0.0168963f $X=9.665 $Y=0.615
+ $X2=0 $Y2=0
cc_840 N_A_1678_395#_c_1223_n N_A_1350_392#_M1032_g 0.00530998f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_841 N_A_1678_395#_c_1226_n N_A_1350_392#_M1032_g 0.00445436f $X=9.722 $Y=1.12
+ $X2=0 $Y2=0
cc_842 N_A_1678_395#_c_1231_n N_A_1350_392#_c_1357_n 0.00748658f $X=9.395
+ $Y=2.445 $X2=0 $Y2=0
cc_843 N_A_1678_395#_c_1232_n N_A_1350_392#_c_1357_n 0.00806887f $X=9.775
+ $Y=1.96 $X2=0 $Y2=0
cc_844 N_A_1678_395#_c_1233_n N_A_1350_392#_c_1357_n 0.00374598f $X=9.48 $Y=1.96
+ $X2=0 $Y2=0
cc_845 N_A_1678_395#_c_1223_n N_A_1350_392#_c_1357_n 0.00340775f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_846 N_A_1678_395#_c_1231_n N_A_1350_392#_c_1358_n 0.00506844f $X=9.395
+ $Y=2.445 $X2=0 $Y2=0
cc_847 N_A_1678_395#_c_1235_n N_A_1350_392#_c_1358_n 0.0087621f $X=9.395
+ $Y=2.675 $X2=0 $Y2=0
cc_848 N_A_1678_395#_c_1223_n N_A_1350_392#_c_1344_n 0.00646442f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_849 N_A_1678_395#_c_1226_n N_A_1350_392#_c_1344_n 0.00210562f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_850 N_A_1678_395#_c_1223_n N_A_1350_392#_c_1360_n 0.00347834f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_851 N_A_1678_395#_c_1231_n N_A_1350_392#_c_1361_n 0.00136199f $X=9.395
+ $Y=2.445 $X2=0 $Y2=0
cc_852 N_A_1678_395#_c_1232_n N_A_1350_392#_c_1361_n 0.00681839f $X=9.775
+ $Y=1.96 $X2=0 $Y2=0
cc_853 N_A_1678_395#_c_1223_n N_A_1350_392#_c_1346_n 2.16647e-19 $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_854 N_A_1678_395#_c_1223_n N_A_1350_392#_c_1347_n 0.00420863f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_855 N_A_1678_395#_c_1226_n N_A_1350_392#_c_1349_n 0.00110652f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_856 N_A_1678_395#_c_1223_n N_A_1350_392#_c_1350_n 0.00382761f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_857 N_A_1678_395#_c_1226_n N_A_1350_392#_c_1350_n 4.03357e-19 $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_858 N_A_1678_395#_c_1228_n N_A_1350_392#_c_1380_n 0.00671391f $X=8.48 $Y=2.39
+ $X2=0 $Y2=0
cc_859 N_A_1678_395#_c_1227_n N_A_1350_392#_c_1368_n 0.00369956f $X=8.48 $Y=2.3
+ $X2=0 $Y2=0
cc_860 N_A_1678_395#_c_1228_n N_A_1350_392#_c_1368_n 0.00436797f $X=8.48 $Y=2.39
+ $X2=0 $Y2=0
cc_861 N_A_1678_395#_c_1220_n N_A_1350_392#_c_1368_n 0.00937113f $X=8.492
+ $Y=1.975 $X2=0 $Y2=0
cc_862 N_A_1678_395#_c_1230_n N_A_1350_392#_c_1368_n 0.00305989f $X=8.492
+ $Y=2.125 $X2=0 $Y2=0
cc_863 N_A_1678_395#_c_1220_n N_A_1350_392#_c_1353_n 0.0106324f $X=8.492
+ $Y=1.975 $X2=0 $Y2=0
cc_864 N_A_1678_395#_c_1230_n N_A_1350_392#_c_1353_n 0.0010085f $X=8.492
+ $Y=2.125 $X2=0 $Y2=0
cc_865 N_A_1678_395#_c_1221_n N_A_1350_392#_c_1353_n 0.0259611f $X=9.5 $Y=1.12
+ $X2=0 $Y2=0
cc_866 N_A_1678_395#_c_1233_n N_A_1350_392#_c_1353_n 0.00291458f $X=9.48 $Y=1.96
+ $X2=0 $Y2=0
cc_867 N_A_1678_395#_c_1224_n N_A_1350_392#_c_1353_n 0.0236067f $X=8.61 $Y=1.12
+ $X2=0 $Y2=0
cc_868 N_A_1678_395#_c_1225_n N_A_1350_392#_c_1353_n 0.00125903f $X=8.61 $Y=1.2
+ $X2=0 $Y2=0
cc_869 N_A_1678_395#_c_1221_n N_A_1350_392#_c_1355_n 0.0111296f $X=9.5 $Y=1.12
+ $X2=0 $Y2=0
cc_870 N_A_1678_395#_c_1232_n N_A_1350_392#_c_1355_n 0.00903277f $X=9.775
+ $Y=1.96 $X2=0 $Y2=0
cc_871 N_A_1678_395#_c_1233_n N_A_1350_392#_c_1355_n 0.0107527f $X=9.48 $Y=1.96
+ $X2=0 $Y2=0
cc_872 N_A_1678_395#_c_1223_n N_A_1350_392#_c_1355_n 0.0237947f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_873 N_A_1678_395#_c_1226_n N_A_1350_392#_c_1355_n 0.00870087f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_874 N_A_1678_395#_c_1221_n N_A_1350_392#_c_1356_n 2.04435e-19 $X=9.5 $Y=1.12
+ $X2=0 $Y2=0
cc_875 N_A_1678_395#_c_1232_n N_A_1350_392#_c_1356_n 0.00306014f $X=9.775
+ $Y=1.96 $X2=0 $Y2=0
cc_876 N_A_1678_395#_c_1233_n N_A_1350_392#_c_1356_n 2.63281e-19 $X=9.48 $Y=1.96
+ $X2=0 $Y2=0
cc_877 N_A_1678_395#_c_1223_n N_A_1350_392#_c_1356_n 0.00218969f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_878 N_A_1678_395#_c_1226_n N_A_1350_392#_c_1356_n 0.00294175f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_879 N_A_1678_395#_c_1231_n N_A_2010_409#_c_1529_n 0.0101593f $X=9.395
+ $Y=2.445 $X2=0 $Y2=0
cc_880 N_A_1678_395#_c_1232_n N_A_2010_409#_c_1529_n 0.0138137f $X=9.775 $Y=1.96
+ $X2=0 $Y2=0
cc_881 N_A_1678_395#_c_1223_n N_A_2010_409#_c_1529_n 0.0176781f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_882 N_A_1678_395#_c_1223_n N_A_2010_409#_c_1518_n 0.0137366f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_883 N_A_1678_395#_c_1223_n N_A_2010_409#_c_1519_n 0.00265607f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_884 N_A_1678_395#_c_1226_n N_A_2010_409#_c_1519_n 0.00237986f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_885 N_A_1678_395#_c_1223_n N_A_2010_409#_c_1521_n 0.00529677f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_886 N_A_1678_395#_c_1232_n N_VPWR_M1008_d 0.00207757f $X=9.775 $Y=1.96 $X2=0
+ $Y2=0
cc_887 N_A_1678_395#_c_1228_n N_VPWR_c_1647_n 0.00418966f $X=8.48 $Y=2.39 $X2=0
+ $Y2=0
cc_888 N_A_1678_395#_c_1230_n N_VPWR_c_1647_n 5.77237e-19 $X=8.492 $Y=2.125
+ $X2=0 $Y2=0
cc_889 N_A_1678_395#_c_1235_n N_VPWR_c_1647_n 0.0193003f $X=9.395 $Y=2.675 $X2=0
+ $Y2=0
cc_890 N_A_1678_395#_c_1232_n N_VPWR_c_1648_n 0.0101135f $X=9.775 $Y=1.96 $X2=0
+ $Y2=0
cc_891 N_A_1678_395#_c_1235_n N_VPWR_c_1648_n 0.0355218f $X=9.395 $Y=2.675 $X2=0
+ $Y2=0
cc_892 N_A_1678_395#_c_1228_n N_VPWR_c_1653_n 0.00519569f $X=8.48 $Y=2.39 $X2=0
+ $Y2=0
cc_893 N_A_1678_395#_c_1235_n N_VPWR_c_1655_n 0.0130061f $X=9.395 $Y=2.675 $X2=0
+ $Y2=0
cc_894 N_A_1678_395#_c_1228_n N_VPWR_c_1640_n 0.0052212f $X=8.48 $Y=2.39 $X2=0
+ $Y2=0
cc_895 N_A_1678_395#_c_1235_n N_VPWR_c_1640_n 0.013771f $X=9.395 $Y=2.675 $X2=0
+ $Y2=0
cc_896 N_A_1678_395#_M1023_g N_VGND_c_2008_n 0.00207012f $X=8.55 $Y=0.615 $X2=0
+ $Y2=0
cc_897 N_A_1678_395#_c_1221_n N_VGND_c_2008_n 0.0139742f $X=9.5 $Y=1.12 $X2=0
+ $Y2=0
cc_898 N_A_1678_395#_c_1222_n N_VGND_c_2008_n 0.00732847f $X=9.665 $Y=0.615
+ $X2=0 $Y2=0
cc_899 N_A_1678_395#_c_1224_n N_VGND_c_2008_n 0.0115305f $X=8.61 $Y=1.12 $X2=0
+ $Y2=0
cc_900 N_A_1678_395#_c_1225_n N_VGND_c_2008_n 0.00115479f $X=8.61 $Y=1.2 $X2=0
+ $Y2=0
cc_901 N_A_1678_395#_c_1222_n N_VGND_c_2009_n 0.0362241f $X=9.665 $Y=0.615 $X2=0
+ $Y2=0
cc_902 N_A_1678_395#_c_1226_n N_VGND_c_2009_n 0.00818535f $X=9.722 $Y=1.12 $X2=0
+ $Y2=0
cc_903 N_A_1678_395#_c_1222_n N_VGND_c_2016_n 0.0127604f $X=9.665 $Y=0.615 $X2=0
+ $Y2=0
cc_904 N_A_1678_395#_M1023_g N_VGND_c_2020_n 0.00551028f $X=8.55 $Y=0.615 $X2=0
+ $Y2=0
cc_905 N_A_1678_395#_M1023_g N_VGND_c_2029_n 0.00534666f $X=8.55 $Y=0.615 $X2=0
+ $Y2=0
cc_906 N_A_1678_395#_c_1222_n N_VGND_c_2029_n 0.011834f $X=9.665 $Y=0.615 $X2=0
+ $Y2=0
cc_907 N_A_1350_392#_c_1363_n N_A_2010_409#_c_1523_n 0.00695913f $X=10.425
+ $Y=1.88 $X2=0 $Y2=0
cc_908 N_A_1350_392#_c_1364_n N_A_2010_409#_c_1523_n 0.0173361f $X=10.425
+ $Y=1.97 $X2=0 $Y2=0
cc_909 N_A_1350_392#_c_1346_n N_A_2010_409#_c_1512_n 0.00125363f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_910 N_A_1350_392#_c_1350_n N_A_2010_409#_c_1512_n 4.19636e-19 $X=10.475
+ $Y=1.335 $X2=0 $Y2=0
cc_911 N_A_1350_392#_c_1346_n N_A_2010_409#_c_1516_n 0.0114635f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_912 N_A_1350_392#_c_1360_n N_A_2010_409#_c_1529_n 0.00194084f $X=9.975
+ $Y=1.88 $X2=0 $Y2=0
cc_913 N_A_1350_392#_c_1361_n N_A_2010_409#_c_1529_n 0.00666311f $X=9.975
+ $Y=1.97 $X2=0 $Y2=0
cc_914 N_A_1350_392#_c_1345_n N_A_2010_409#_c_1529_n 0.00471727f $X=10.335
+ $Y=1.63 $X2=0 $Y2=0
cc_915 N_A_1350_392#_c_1363_n N_A_2010_409#_c_1529_n 0.0049772f $X=10.425
+ $Y=1.88 $X2=0 $Y2=0
cc_916 N_A_1350_392#_c_1364_n N_A_2010_409#_c_1529_n 0.0151283f $X=10.425
+ $Y=1.97 $X2=0 $Y2=0
cc_917 N_A_1350_392#_c_1348_n N_A_2010_409#_c_1529_n 0.00143923f $X=10.425
+ $Y=1.63 $X2=0 $Y2=0
cc_918 N_A_1350_392#_c_1346_n N_A_2010_409#_c_1517_n 0.00840659f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_919 N_A_1350_392#_c_1348_n N_A_2010_409#_c_1517_n 0.00857014f $X=10.425
+ $Y=1.63 $X2=0 $Y2=0
cc_920 N_A_1350_392#_c_1350_n N_A_2010_409#_c_1517_n 0.00194299f $X=10.475
+ $Y=1.335 $X2=0 $Y2=0
cc_921 N_A_1350_392#_c_1345_n N_A_2010_409#_c_1518_n 0.00614927f $X=10.335
+ $Y=1.63 $X2=0 $Y2=0
cc_922 N_A_1350_392#_c_1346_n N_A_2010_409#_c_1518_n 0.00148617f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_923 N_A_1350_392#_c_1348_n N_A_2010_409#_c_1518_n 6.95643e-19 $X=10.425
+ $Y=1.63 $X2=0 $Y2=0
cc_924 N_A_1350_392#_c_1349_n N_A_2010_409#_c_1519_n 0.0127757f $X=10.475
+ $Y=1.185 $X2=0 $Y2=0
cc_925 N_A_1350_392#_c_1350_n N_A_2010_409#_c_1519_n 0.00490997f $X=10.475
+ $Y=1.335 $X2=0 $Y2=0
cc_926 N_A_1350_392#_c_1346_n N_A_2010_409#_c_1521_n 0.0026095f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_927 N_A_1350_392#_c_1350_n N_A_2010_409#_c_1521_n 0.00200729f $X=10.475
+ $Y=1.335 $X2=0 $Y2=0
cc_928 N_A_1350_392#_c_1368_n N_VPWR_c_1647_n 0.0017733f $X=8.325 $Y=2.475 $X2=0
+ $Y2=0
cc_929 N_A_1350_392#_c_1358_n N_VPWR_c_1648_n 0.00436524f $X=9.47 $Y=2.39 $X2=0
+ $Y2=0
cc_930 N_A_1350_392#_c_1361_n N_VPWR_c_1648_n 0.00225694f $X=9.975 $Y=1.97 $X2=0
+ $Y2=0
cc_931 N_A_1350_392#_c_1364_n N_VPWR_c_1649_n 0.00658928f $X=10.425 $Y=1.97
+ $X2=0 $Y2=0
cc_932 N_A_1350_392#_c_1351_n N_VPWR_c_1653_n 0.00505902f $X=7.245 $Y=2.475
+ $X2=0 $Y2=0
cc_933 N_A_1350_392#_c_1380_n N_VPWR_c_1653_n 0.0236614f $X=8.24 $Y=2.64 $X2=0
+ $Y2=0
cc_934 N_A_1350_392#_c_1358_n N_VPWR_c_1655_n 0.0044306f $X=9.47 $Y=2.39 $X2=0
+ $Y2=0
cc_935 N_A_1350_392#_c_1361_n N_VPWR_c_1657_n 0.00522765f $X=9.975 $Y=1.97 $X2=0
+ $Y2=0
cc_936 N_A_1350_392#_c_1364_n N_VPWR_c_1657_n 0.00510653f $X=10.425 $Y=1.97
+ $X2=0 $Y2=0
cc_937 N_A_1350_392#_c_1358_n N_VPWR_c_1640_n 0.0052212f $X=9.47 $Y=2.39 $X2=0
+ $Y2=0
cc_938 N_A_1350_392#_c_1361_n N_VPWR_c_1640_n 0.0052212f $X=9.975 $Y=1.97 $X2=0
+ $Y2=0
cc_939 N_A_1350_392#_c_1364_n N_VPWR_c_1640_n 0.0052212f $X=10.425 $Y=1.97 $X2=0
+ $Y2=0
cc_940 N_A_1350_392#_c_1351_n N_VPWR_c_1640_n 0.00669727f $X=7.245 $Y=2.475
+ $X2=0 $Y2=0
cc_941 N_A_1350_392#_c_1380_n N_VPWR_c_1640_n 0.0343965f $X=8.24 $Y=2.64 $X2=0
+ $Y2=0
cc_942 N_A_1350_392#_c_1380_n A_1627_493# 0.00324022f $X=8.24 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_943 N_A_1350_392#_M1032_g N_VGND_c_2009_n 0.00460851f $X=9.45 $Y=0.615 $X2=0
+ $Y2=0
cc_944 N_A_1350_392#_c_1345_n N_VGND_c_2009_n 0.00151024f $X=10.335 $Y=1.63
+ $X2=0 $Y2=0
cc_945 N_A_1350_392#_c_1349_n N_VGND_c_2009_n 0.0197658f $X=10.475 $Y=1.185
+ $X2=0 $Y2=0
cc_946 N_A_1350_392#_c_1350_n N_VGND_c_2009_n 8.25701e-19 $X=10.475 $Y=1.335
+ $X2=0 $Y2=0
cc_947 N_A_1350_392#_c_1349_n N_VGND_c_2010_n 0.00422452f $X=10.475 $Y=1.185
+ $X2=0 $Y2=0
cc_948 N_A_1350_392#_M1032_g N_VGND_c_2016_n 0.00527282f $X=9.45 $Y=0.615 $X2=0
+ $Y2=0
cc_949 N_A_1350_392#_c_1349_n N_VGND_c_2021_n 0.00434272f $X=10.475 $Y=1.185
+ $X2=0 $Y2=0
cc_950 N_A_1350_392#_M1032_g N_VGND_c_2029_n 0.00534666f $X=9.45 $Y=0.615 $X2=0
+ $Y2=0
cc_951 N_A_1350_392#_c_1349_n N_VGND_c_2029_n 0.00830058f $X=10.475 $Y=1.185
+ $X2=0 $Y2=0
cc_952 N_A_2010_409#_c_1529_n N_VPWR_c_1648_n 0.028739f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_953 N_A_2010_409#_c_1523_n N_VPWR_c_1649_n 0.0157125f $X=10.93 $Y=1.765 $X2=0
+ $Y2=0
cc_954 N_A_2010_409#_c_1524_n N_VPWR_c_1649_n 5.87659e-19 $X=11.425 $Y=1.765
+ $X2=0 $Y2=0
cc_955 N_A_2010_409#_c_1529_n N_VPWR_c_1649_n 0.0332253f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_956 N_A_2010_409#_c_1517_n N_VPWR_c_1649_n 0.00110837f $X=10.56 $Y=1.545
+ $X2=0 $Y2=0
cc_957 N_A_2010_409#_c_1521_n N_VPWR_c_1649_n 0.0137726f $X=10.725 $Y=1.465
+ $X2=0 $Y2=0
cc_958 N_A_2010_409#_c_1524_n N_VPWR_c_1650_n 0.00634007f $X=11.425 $Y=1.765
+ $X2=0 $Y2=0
cc_959 N_A_2010_409#_c_1526_n N_VPWR_c_1650_n 0.00634007f $X=12.35 $Y=1.765
+ $X2=0 $Y2=0
cc_960 N_A_2010_409#_c_1527_n N_VPWR_c_1652_n 0.0235387f $X=12.8 $Y=1.765 $X2=0
+ $Y2=0
cc_961 N_A_2010_409#_c_1522_n N_VPWR_c_1652_n 6.01683e-19 $X=12.8 $Y=1.532 $X2=0
+ $Y2=0
cc_962 N_A_2010_409#_c_1529_n N_VPWR_c_1657_n 0.00845353f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_963 N_A_2010_409#_c_1523_n N_VPWR_c_1663_n 0.00429299f $X=10.93 $Y=1.765
+ $X2=0 $Y2=0
cc_964 N_A_2010_409#_c_1524_n N_VPWR_c_1663_n 0.00445602f $X=11.425 $Y=1.765
+ $X2=0 $Y2=0
cc_965 N_A_2010_409#_c_1526_n N_VPWR_c_1664_n 0.00445602f $X=12.35 $Y=1.765
+ $X2=0 $Y2=0
cc_966 N_A_2010_409#_c_1527_n N_VPWR_c_1664_n 0.00445602f $X=12.8 $Y=1.765 $X2=0
+ $Y2=0
cc_967 N_A_2010_409#_c_1523_n N_VPWR_c_1640_n 0.00848138f $X=10.93 $Y=1.765
+ $X2=0 $Y2=0
cc_968 N_A_2010_409#_c_1524_n N_VPWR_c_1640_n 0.00862136f $X=11.425 $Y=1.765
+ $X2=0 $Y2=0
cc_969 N_A_2010_409#_c_1526_n N_VPWR_c_1640_n 0.00861719f $X=12.35 $Y=1.765
+ $X2=0 $Y2=0
cc_970 N_A_2010_409#_c_1527_n N_VPWR_c_1640_n 0.00860781f $X=12.8 $Y=1.765 $X2=0
+ $Y2=0
cc_971 N_A_2010_409#_c_1529_n N_VPWR_c_1640_n 0.00872066f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_972 N_A_2010_409#_c_1523_n N_Q_c_1939_n 4.36646e-19 $X=10.93 $Y=1.765 $X2=0
+ $Y2=0
cc_973 N_A_2010_409#_c_1524_n N_Q_c_1939_n 0.0165329f $X=11.425 $Y=1.765 $X2=0
+ $Y2=0
cc_974 N_A_2010_409#_c_1524_n N_Q_c_1940_n 0.0139279f $X=11.425 $Y=1.765 $X2=0
+ $Y2=0
cc_975 N_A_2010_409#_c_1512_n N_Q_c_1940_n 0.018687f $X=11.575 $Y=1.465 $X2=0
+ $Y2=0
cc_976 N_A_2010_409#_c_1526_n N_Q_c_1940_n 0.0152854f $X=12.35 $Y=1.765 $X2=0
+ $Y2=0
cc_977 N_A_2010_409#_c_1520_n N_Q_c_1940_n 0.0651475f $X=12.075 $Y=1.465 $X2=0
+ $Y2=0
cc_978 N_A_2010_409#_c_1522_n N_Q_c_1940_n 4.77499e-19 $X=12.8 $Y=1.532 $X2=0
+ $Y2=0
cc_979 N_A_2010_409#_c_1523_n N_Q_c_1941_n 7.16209e-19 $X=10.93 $Y=1.765 $X2=0
+ $Y2=0
cc_980 N_A_2010_409#_c_1509_n N_Q_c_1941_n 0.00632181f $X=11.23 $Y=1.555 $X2=0
+ $Y2=0
cc_981 N_A_2010_409#_c_1524_n N_Q_c_1941_n 9.16146e-19 $X=11.425 $Y=1.765 $X2=0
+ $Y2=0
cc_982 N_A_2010_409#_c_1512_n N_Q_c_1941_n 4.41065e-19 $X=11.575 $Y=1.465 $X2=0
+ $Y2=0
cc_983 N_A_2010_409#_c_1529_n N_Q_c_1941_n 0.00261306f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_984 N_A_2010_409#_c_1520_n N_Q_c_1941_n 0.0277245f $X=12.075 $Y=1.465 $X2=0
+ $Y2=0
cc_985 N_A_2010_409#_M1003_g N_Q_c_1932_n 2.01997e-19 $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_986 N_A_2010_409#_c_1511_n N_Q_c_1932_n 0.00454265f $X=11.95 $Y=1.465 $X2=0
+ $Y2=0
cc_987 N_A_2010_409#_c_1520_n N_Q_c_1932_n 0.0265674f $X=12.075 $Y=1.465 $X2=0
+ $Y2=0
cc_988 N_A_2010_409#_M1003_g N_Q_c_1933_n 3.0578e-19 $X=11.5 $Y=0.74 $X2=0 $Y2=0
cc_989 N_A_2010_409#_M1024_g N_Q_c_1933_n 2.92386e-19 $X=12.025 $Y=0.74 $X2=0
+ $Y2=0
cc_990 N_A_2010_409#_M1024_g N_Q_c_1934_n 0.0154071f $X=12.025 $Y=0.74 $X2=0
+ $Y2=0
cc_991 N_A_2010_409#_M1033_g N_Q_c_1934_n 0.0148564f $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_992 N_A_2010_409#_c_1520_n N_Q_c_1934_n 0.0248822f $X=12.075 $Y=1.465 $X2=0
+ $Y2=0
cc_993 N_A_2010_409#_c_1522_n N_Q_c_1934_n 0.00819925f $X=12.8 $Y=1.532 $X2=0
+ $Y2=0
cc_994 N_A_2010_409#_c_1526_n N_Q_c_1942_n 0.0165744f $X=12.35 $Y=1.765 $X2=0
+ $Y2=0
cc_995 N_A_2010_409#_c_1527_n N_Q_c_1942_n 0.011071f $X=12.8 $Y=1.765 $X2=0
+ $Y2=0
cc_996 N_A_2010_409#_M1024_g N_Q_c_1935_n 5.92753e-19 $X=12.025 $Y=0.74 $X2=0
+ $Y2=0
cc_997 N_A_2010_409#_M1033_g N_Q_c_1935_n 0.00800161f $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_998 N_A_2010_409#_M1038_g N_Q_c_1935_n 3.97481e-19 $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_999 N_A_2010_409#_M1024_g N_Q_c_1936_n 6.59139e-19 $X=12.025 $Y=0.74 $X2=0
+ $Y2=0
cc_1000 N_A_2010_409#_M1033_g N_Q_c_1936_n 0.00385048f $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_1001 N_A_2010_409#_M1038_g N_Q_c_1936_n 0.00355386f $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1002 N_A_2010_409#_M1033_g N_Q_c_1937_n 7.39274e-19 $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_1003 N_A_2010_409#_M1038_g N_Q_c_1937_n 6.05444e-19 $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1004 N_A_2010_409#_c_1526_n Q 0.00265569f $X=12.35 $Y=1.765 $X2=0 $Y2=0
cc_1005 N_A_2010_409#_M1033_g Q 0.0055056f $X=12.525 $Y=0.74 $X2=0 $Y2=0
cc_1006 N_A_2010_409#_c_1527_n Q 0.0163525f $X=12.8 $Y=1.765 $X2=0 $Y2=0
cc_1007 N_A_2010_409#_M1038_g Q 0.0162652f $X=12.955 $Y=0.74 $X2=0 $Y2=0
cc_1008 N_A_2010_409#_c_1520_n Q 0.0167026f $X=12.075 $Y=1.465 $X2=0 $Y2=0
cc_1009 N_A_2010_409#_c_1522_n Q 0.0439249f $X=12.8 $Y=1.532 $X2=0 $Y2=0
cc_1010 N_A_2010_409#_c_1517_n N_VGND_c_2009_n 0.00116291f $X=10.56 $Y=1.545
+ $X2=0 $Y2=0
cc_1011 N_A_2010_409#_c_1518_n N_VGND_c_2009_n 0.0146779f $X=10.365 $Y=1.545
+ $X2=0 $Y2=0
cc_1012 N_A_2010_409#_c_1519_n N_VGND_c_2009_n 0.0308054f $X=10.725 $Y=0.515
+ $X2=0 $Y2=0
cc_1013 N_A_2010_409#_c_1509_n N_VGND_c_2010_n 5.70705e-19 $X=11.23 $Y=1.555
+ $X2=0 $Y2=0
cc_1014 N_A_2010_409#_M1003_g N_VGND_c_2010_n 0.00531367f $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_1015 N_A_2010_409#_c_1512_n N_VGND_c_2010_n 0.00442734f $X=11.575 $Y=1.465
+ $X2=0 $Y2=0
cc_1016 N_A_2010_409#_c_1519_n N_VGND_c_2010_n 0.0520772f $X=10.725 $Y=0.515
+ $X2=0 $Y2=0
cc_1017 N_A_2010_409#_c_1520_n N_VGND_c_2010_n 0.0247375f $X=12.075 $Y=1.465
+ $X2=0 $Y2=0
cc_1018 N_A_2010_409#_M1003_g N_VGND_c_2011_n 4.65028e-19 $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_1019 N_A_2010_409#_M1024_g N_VGND_c_2011_n 0.00807752f $X=12.025 $Y=0.74
+ $X2=0 $Y2=0
cc_1020 N_A_2010_409#_M1033_g N_VGND_c_2011_n 0.00355746f $X=12.525 $Y=0.74
+ $X2=0 $Y2=0
cc_1021 N_A_2010_409#_M1033_g N_VGND_c_2013_n 5.9507e-19 $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_1022 N_A_2010_409#_M1038_g N_VGND_c_2013_n 0.0138049f $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1023 N_A_2010_409#_c_1519_n N_VGND_c_2021_n 0.0145639f $X=10.725 $Y=0.515
+ $X2=0 $Y2=0
cc_1024 N_A_2010_409#_M1003_g N_VGND_c_2022_n 0.00461464f $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_1025 N_A_2010_409#_M1024_g N_VGND_c_2022_n 0.00398535f $X=12.025 $Y=0.74
+ $X2=0 $Y2=0
cc_1026 N_A_2010_409#_M1033_g N_VGND_c_2023_n 0.00434272f $X=12.525 $Y=0.74
+ $X2=0 $Y2=0
cc_1027 N_A_2010_409#_M1038_g N_VGND_c_2023_n 0.00383152f $X=12.955 $Y=0.74
+ $X2=0 $Y2=0
cc_1028 N_A_2010_409#_M1003_g N_VGND_c_2029_n 0.00913308f $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_1029 N_A_2010_409#_M1024_g N_VGND_c_2029_n 0.00788407f $X=12.025 $Y=0.74
+ $X2=0 $Y2=0
cc_1030 N_A_2010_409#_M1033_g N_VGND_c_2029_n 0.00820718f $X=12.525 $Y=0.74
+ $X2=0 $Y2=0
cc_1031 N_A_2010_409#_M1038_g N_VGND_c_2029_n 0.0075754f $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1032 N_A_2010_409#_c_1519_n N_VGND_c_2029_n 0.0119984f $X=10.725 $Y=0.515
+ $X2=0 $Y2=0
cc_1033 N_VPWR_M1004_d N_A_37_78#_c_1813_n 0.00501542f $X=2.02 $Y=1.83 $X2=0
+ $Y2=0
cc_1034 N_VPWR_c_1644_n N_A_37_78#_c_1813_n 0.0162734f $X=2.17 $Y=2.785 $X2=0
+ $Y2=0
cc_1035 N_VPWR_c_1640_n N_A_37_78#_c_1813_n 0.0238036f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1036 N_VPWR_c_1642_n N_A_37_78#_c_1816_n 0.0310355f $X=0.275 $Y=2.75 $X2=0
+ $Y2=0
cc_1037 N_VPWR_c_1643_n N_A_37_78#_c_1816_n 0.0222518f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_1038 N_VPWR_c_1659_n N_A_37_78#_c_1816_n 0.0144812f $X=1.09 $Y=3.33 $X2=0
+ $Y2=0
cc_1039 N_VPWR_c_1640_n N_A_37_78#_c_1816_n 0.0119834f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1040 N_VPWR_c_1643_n N_A_37_78#_c_1817_n 0.0193352f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_1041 N_VPWR_c_1640_n N_A_37_78#_c_1817_n 0.0125344f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1042 N_VPWR_c_1640_n N_A_37_78#_c_1818_n 0.0170528f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1043 N_VPWR_c_1661_n N_A_37_78#_c_1819_n 0.007532f $X=4.4 $Y=3.33 $X2=0 $Y2=0
cc_1044 N_VPWR_c_1640_n N_A_37_78#_c_1819_n 0.00909433f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1045 N_VPWR_c_1649_n N_Q_c_1939_n 0.0366244f $X=10.7 $Y=2.19 $X2=0 $Y2=0
cc_1046 N_VPWR_c_1650_n N_Q_c_1939_n 0.0324053f $X=12.12 $Y=2.305 $X2=0 $Y2=0
cc_1047 N_VPWR_c_1663_n N_Q_c_1939_n 0.0145938f $X=11.535 $Y=3.33 $X2=0 $Y2=0
cc_1048 N_VPWR_c_1640_n N_Q_c_1939_n 0.0120466f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1049 N_VPWR_M1013_s N_Q_c_1940_n 0.00998974f $X=11.5 $Y=1.84 $X2=0 $Y2=0
cc_1050 N_VPWR_c_1650_n N_Q_c_1940_n 0.053778f $X=12.12 $Y=2.305 $X2=0 $Y2=0
cc_1051 N_VPWR_c_1650_n N_Q_c_1942_n 0.0324053f $X=12.12 $Y=2.305 $X2=0 $Y2=0
cc_1052 N_VPWR_c_1652_n N_Q_c_1942_n 0.0386506f $X=13.075 $Y=2.115 $X2=0 $Y2=0
cc_1053 N_VPWR_c_1664_n N_Q_c_1942_n 0.014552f $X=12.91 $Y=3.33 $X2=0 $Y2=0
cc_1054 N_VPWR_c_1640_n N_Q_c_1942_n 0.0119791f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1055 N_VPWR_c_1652_n Q 0.0285893f $X=13.075 $Y=2.115 $X2=0 $Y2=0
cc_1056 N_A_37_78#_c_1805_n A_124_78# 0.00236678f $X=0.685 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_1057 N_A_37_78#_c_1805_n N_VGND_c_2006_n 0.00131521f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_1058 N_A_37_78#_c_1811_n N_VGND_c_2006_n 0.00434714f $X=0.33 $Y=0.6 $X2=0
+ $Y2=0
cc_1059 N_A_37_78#_c_1805_n N_VGND_c_2014_n 0.00520932f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_1060 N_A_37_78#_c_1811_n N_VGND_c_2014_n 0.0131067f $X=0.33 $Y=0.6 $X2=0
+ $Y2=0
cc_1061 N_A_37_78#_c_1805_n N_VGND_c_2029_n 0.0102476f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_1062 N_A_37_78#_c_1811_n N_VGND_c_2029_n 0.0117869f $X=0.33 $Y=0.6 $X2=0
+ $Y2=0
cc_1063 N_Q_c_1934_n N_VGND_M1024_d 0.00253871f $X=12.575 $Y=1.005 $X2=0 $Y2=0
cc_1064 N_Q_c_1932_n N_VGND_c_2010_n 0.00156718f $X=11.752 $Y=0.88 $X2=0 $Y2=0
cc_1065 N_Q_c_1933_n N_VGND_c_2010_n 3.09414e-19 $X=11.76 $Y=0.53 $X2=0 $Y2=0
cc_1066 N_Q_c_1933_n N_VGND_c_2011_n 0.0130802f $X=11.76 $Y=0.53 $X2=0 $Y2=0
cc_1067 N_Q_c_1934_n N_VGND_c_2011_n 0.0211572f $X=12.575 $Y=1.005 $X2=0 $Y2=0
cc_1068 N_Q_c_1935_n N_VGND_c_2011_n 0.0137341f $X=12.74 $Y=0.515 $X2=0 $Y2=0
cc_1069 N_Q_c_1935_n N_VGND_c_2013_n 0.0197239f $X=12.74 $Y=0.515 $X2=0 $Y2=0
cc_1070 Q N_VGND_c_2013_n 0.0250286f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_1071 N_Q_c_1933_n N_VGND_c_2022_n 0.0131726f $X=11.76 $Y=0.53 $X2=0 $Y2=0
cc_1072 N_Q_c_1935_n N_VGND_c_2023_n 0.0109942f $X=12.74 $Y=0.515 $X2=0 $Y2=0
cc_1073 N_Q_c_1933_n N_VGND_c_2029_n 0.0114552f $X=11.76 $Y=0.53 $X2=0 $Y2=0
cc_1074 N_Q_c_1935_n N_VGND_c_2029_n 0.00904371f $X=12.74 $Y=0.515 $X2=0 $Y2=0
