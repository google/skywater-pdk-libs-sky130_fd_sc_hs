* File: sky130_fd_sc_hs__o221a_4.pex.spice
* Created: Thu Aug 27 20:59:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O221A_4%C1 3 5 7 10 12 14 15 16 24
c47 10 0 1.44963e-19 $X=0.925 $Y=0.945
r48 24 25 3.94005 $w=3.67e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.652
+ $X2=0.955 $Y2=1.652
r49 22 24 26.267 $w=3.67e-07 $l=2e-07 $layer=POLY_cond $X=0.725 $Y=1.652
+ $X2=0.925 $Y2=1.652
r50 20 22 28.8937 $w=3.67e-07 $l=2.2e-07 $layer=POLY_cond $X=0.505 $Y=1.652
+ $X2=0.725 $Y2=1.652
r51 19 20 1.31335 $w=3.67e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.652
+ $X2=0.505 $Y2=1.652
r52 16 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.61 $X2=0.725 $Y2=1.61
r53 15 16 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.612
+ $X2=0.72 $Y2=1.612
r54 12 25 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.86
+ $X2=0.955 $Y2=1.652
r55 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.86
+ $X2=0.955 $Y2=2.435
r56 8 24 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.445
+ $X2=0.925 $Y2=1.652
r57 8 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.925 $Y=1.445
+ $X2=0.925 $Y2=0.945
r58 5 20 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.86
+ $X2=0.505 $Y2=1.652
r59 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.86
+ $X2=0.505 $Y2=2.435
r60 1 19 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.445
+ $X2=0.495 $Y2=1.652
r61 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.495 $Y=1.445 $X2=0.495
+ $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%B2 3 5 7 10 12 14 15 16 24
c52 24 0 8.30843e-20 $X=2.355 $Y=1.652
c53 16 0 1.5371e-19 $X=2.64 $Y=1.665
c54 3 0 1.70191e-19 $X=1.89 $Y=0.945
r55 22 24 9.56349 $w=3.78e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=1.652
+ $X2=2.355 $Y2=1.652
r56 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.61 $X2=2.28 $Y2=1.61
r57 20 22 47.8175 $w=3.78e-07 $l=3.75e-07 $layer=POLY_cond $X=1.905 $Y=1.652
+ $X2=2.28 $Y2=1.652
r58 19 20 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=1.89 $Y=1.652
+ $X2=1.905 $Y2=1.652
r59 16 23 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=2.64 $Y=1.612
+ $X2=2.28 $Y2=1.612
r60 15 23 4.12815 $w=3.33e-07 $l=1.2e-07 $layer=LI1_cond $X=2.16 $Y=1.612
+ $X2=2.28 $Y2=1.612
r61 12 24 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.355 $Y=1.86
+ $X2=2.355 $Y2=1.652
r62 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.355 $Y=1.86
+ $X2=2.355 $Y2=2.435
r63 8 24 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.355 $Y=1.445
+ $X2=2.355 $Y2=1.652
r64 8 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.355 $Y=1.445
+ $X2=2.355 $Y2=0.945
r65 5 20 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.86
+ $X2=1.905 $Y2=1.652
r66 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.86
+ $X2=1.905 $Y2=2.435
r67 1 19 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.89 $Y=1.445
+ $X2=1.89 $Y2=1.652
r68 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.89 $Y=1.445 $X2=1.89
+ $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%B1 1 2 3 5 9 10 11 14 17 18 20 24 26 27 28
+ 29 36 37
c90 37 0 1.5371e-19 $X=3.3 $Y=1.61
c91 29 0 8.30843e-20 $X=4.08 $Y=1.665
r92 34 37 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.27 $Y=1.61 $X2=3.3
+ $Y2=1.61
r93 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.61
+ $X2=3.105 $Y2=1.61
r94 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.61 $X2=3.27 $Y2=1.61
r95 28 29 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.612
+ $X2=4.08 $Y2=1.612
r96 28 35 11.3524 $w=3.33e-07 $l=3.3e-07 $layer=LI1_cond $X=3.6 $Y=1.612
+ $X2=3.27 $Y2=1.612
r97 27 35 5.16019 $w=3.33e-07 $l=1.5e-07 $layer=LI1_cond $X=3.12 $Y=1.612
+ $X2=3.27 $Y2=1.612
r98 24 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.445
+ $X2=3.3 $Y2=1.61
r99 23 24 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=3.3 $Y=0.255
+ $X2=3.3 $Y2=1.445
r100 22 26 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.895 $Y=1.52
+ $X2=2.805 $Y2=1.52
r101 22 36 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.895 $Y=1.52
+ $X2=3.105 $Y2=1.52
r102 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.805 $Y=1.86
+ $X2=2.805 $Y2=2.435
r103 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.805 $Y=1.77
+ $X2=2.805 $Y2=1.86
r104 16 26 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.805 $Y=1.595
+ $X2=2.805 $Y2=1.52
r105 16 17 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.805 $Y=1.595
+ $X2=2.805 $Y2=1.77
r106 12 26 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.79 $Y=1.445
+ $X2=2.805 $Y2=1.52
r107 12 14 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.79 $Y=1.445
+ $X2=2.79 $Y2=0.945
r108 10 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.225 $Y=0.18
+ $X2=3.3 $Y2=0.255
r109 10 11 884.521 $w=1.5e-07 $l=1.725e-06 $layer=POLY_cond $X=3.225 $Y=0.18
+ $X2=1.5 $Y2=0.18
r110 9 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.425 $Y=0.945
+ $X2=1.425 $Y2=1.34
r111 6 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.425 $Y=0.255
+ $X2=1.5 $Y2=0.18
r112 6 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.425 $Y=0.255
+ $X2=1.425 $Y2=0.945
r113 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.41 $Y=1.86
+ $X2=1.41 $Y2=2.435
r114 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.41 $Y=1.77 $X2=1.41
+ $Y2=1.86
r115 1 25 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.41 $Y=1.43 $X2=1.41
+ $Y2=1.34
r116 1 2 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.41 $Y=1.43 $X2=1.41
+ $Y2=1.77
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%A2 1 3 6 10 12 14 15 22
c44 15 0 1.7872e-19 $X=4.56 $Y=1.665
c45 10 0 3.38411e-20 $X=4.675 $Y=0.915
c46 6 0 6.92713e-20 $X=4.245 $Y=0.915
r47 22 23 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=4.675 $Y=1.652
+ $X2=4.69 $Y2=1.652
r48 20 22 18.9404 $w=3.69e-07 $l=1.45e-07 $layer=POLY_cond $X=4.53 $Y=1.652
+ $X2=4.675 $Y2=1.652
r49 18 20 37.2276 $w=3.69e-07 $l=2.85e-07 $layer=POLY_cond $X=4.245 $Y=1.652
+ $X2=4.53 $Y2=1.652
r50 17 18 3.9187 $w=3.69e-07 $l=3e-08 $layer=POLY_cond $X=4.215 $Y=1.652
+ $X2=4.245 $Y2=1.652
r51 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.61 $X2=4.53 $Y2=1.61
r52 12 23 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.69 $Y=1.86
+ $X2=4.69 $Y2=1.652
r53 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.69 $Y=1.86
+ $X2=4.69 $Y2=2.435
r54 8 22 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.675 $Y=1.445
+ $X2=4.675 $Y2=1.652
r55 8 10 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.675 $Y=1.445
+ $X2=4.675 $Y2=0.915
r56 4 18 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.245 $Y=1.445
+ $X2=4.245 $Y2=1.652
r57 4 6 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.245 $Y=1.445
+ $X2=4.245 $Y2=0.915
r58 1 17 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.215 $Y=1.86
+ $X2=4.215 $Y2=1.652
r59 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.215 $Y=1.86
+ $X2=4.215 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%A1 2 3 5 9 10 11 15 16 18 20 21 25
c74 25 0 4.13126e-20 $X=5.155 $Y=1.515
c75 20 0 1.48608e-19 $X=3.767 $Y=1.46
c76 9 0 2.67289e-19 $X=3.81 $Y=0.915
c77 2 0 1.70982e-19 $X=3.74 $Y=1.77
r78 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.515 $X2=5.155 $Y2=1.515
r79 21 25 4.37637 $w=3.93e-07 $l=1.5e-07 $layer=LI1_cond $X=5.122 $Y=1.665
+ $X2=5.122 $Y2=1.515
r80 19 20 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.767 $Y=1.31
+ $X2=3.767 $Y2=1.46
r81 16 24 70.0964 $w=2.77e-07 $l=3.62077e-07 $layer=POLY_cond $X=5.19 $Y=1.86
+ $X2=5.155 $Y2=1.515
r82 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.19 $Y=1.86
+ $X2=5.19 $Y2=2.435
r83 13 24 38.7751 $w=2.77e-07 $l=1.88348e-07 $layer=POLY_cond $X=5.105 $Y=1.35
+ $X2=5.155 $Y2=1.515
r84 13 15 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.105 $Y=1.35
+ $X2=5.105 $Y2=0.915
r85 12 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.105 $Y=0.255
+ $X2=5.105 $Y2=0.915
r86 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.03 $Y=0.18
+ $X2=5.105 $Y2=0.255
r87 10 11 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=5.03 $Y=0.18
+ $X2=3.885 $Y2=0.18
r88 9 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.81 $Y=0.915
+ $X2=3.81 $Y2=1.31
r89 6 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.81 $Y=0.255
+ $X2=3.885 $Y2=0.18
r90 6 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.81 $Y=0.255 $X2=3.81
+ $Y2=0.915
r91 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.74 $Y=1.86 $X2=3.74
+ $Y2=2.435
r92 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.74 $Y=1.77 $X2=3.74
+ $Y2=1.86
r93 2 20 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=3.74 $Y=1.77 $X2=3.74
+ $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%A_114_125# 1 2 3 4 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 32 33 35 36 38 42 46 48 49 51 52 53 56 60 63 64 69 77 79
c182 64 0 1.22796e-19 $X=5.66 $Y=1.515
c183 56 0 1.40871e-19 $X=4.3 $Y=2.035
c184 42 0 1.44963e-19 $X=0.71 $Y=0.77
c185 19 0 1.46284e-19 $X=6.115 $Y=1.35
c186 16 0 1.65088e-19 $X=5.695 $Y=1.765
r187 86 87 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=6.67 $Y=1.557
+ $X2=6.685 $Y2=1.557
r188 83 84 13.7154 $w=3.69e-07 $l=1.05e-07 $layer=POLY_cond $X=6.115 $Y=1.557
+ $X2=6.22 $Y2=1.557
r189 80 81 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=5.68 $Y=1.557
+ $X2=5.695 $Y2=1.557
r190 73 75 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.73 $Y=2.035
+ $X2=1.145 $Y2=2.035
r191 70 86 28.7371 $w=3.69e-07 $l=2.2e-07 $layer=POLY_cond $X=6.45 $Y=1.557
+ $X2=6.67 $Y2=1.557
r192 70 84 30.0434 $w=3.69e-07 $l=2.3e-07 $layer=POLY_cond $X=6.45 $Y=1.557
+ $X2=6.22 $Y2=1.557
r193 69 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.515 $X2=6.45 $Y2=1.515
r194 67 83 45.065 $w=3.69e-07 $l=3.45e-07 $layer=POLY_cond $X=5.77 $Y=1.557
+ $X2=6.115 $Y2=1.557
r195 67 81 9.79675 $w=3.69e-07 $l=7.5e-08 $layer=POLY_cond $X=5.77 $Y=1.557
+ $X2=5.695 $Y2=1.557
r196 66 69 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.77 $Y=1.515
+ $X2=6.45 $Y2=1.515
r197 66 67 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.77
+ $Y=1.515 $X2=5.77 $Y2=1.515
r198 64 66 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.66 $Y=1.515
+ $X2=5.77 $Y2=1.515
r199 62 64 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.575 $Y=1.68
+ $X2=5.66 $Y2=1.515
r200 62 63 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.575 $Y=1.68
+ $X2=5.575 $Y2=1.95
r201 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=2.035
+ $X2=4.465 $Y2=2.035
r202 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.49 $Y=2.035
+ $X2=5.575 $Y2=1.95
r203 60 61 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.49 $Y=2.035
+ $X2=4.63 $Y2=2.035
r204 57 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=2.035
+ $X2=2.13 $Y2=2.035
r205 56 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=2.035
+ $X2=4.465 $Y2=2.035
r206 56 57 136.027 $w=1.68e-07 $l=2.085e-06 $layer=LI1_cond $X=4.3 $Y=2.035
+ $X2=2.215 $Y2=2.035
r207 53 75 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.035
+ $X2=1.145 $Y2=2.035
r208 52 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.13 $Y2=2.035
r209 52 53 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=1.23 $Y2=2.035
r210 51 75 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.95
+ $X2=1.145 $Y2=2.035
r211 50 51 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.145 $Y=1.275
+ $X2=1.145 $Y2=1.95
r212 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=1.19
+ $X2=1.145 $Y2=1.275
r213 48 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.06 $Y=1.19
+ $X2=0.795 $Y2=1.19
r214 46 73 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=0.73 $Y=2.79
+ $X2=0.73 $Y2=2.12
r215 40 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.67 $Y=1.105
+ $X2=0.795 $Y2=1.19
r216 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.67 $Y=1.105
+ $X2=0.67 $Y2=0.77
r217 36 38 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.175 $Y=1.765
+ $X2=7.175 $Y2=2.4
r218 33 35 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.115 $Y=1.35
+ $X2=7.115 $Y2=0.865
r219 32 87 13.0285 $w=3.69e-07 $l=1.04283e-07 $layer=POLY_cond $X=6.76 $Y=1.487
+ $X2=6.685 $Y2=1.557
r220 31 36 68.0294 $w=2.09e-07 $l=2.89271e-07 $layer=POLY_cond $X=7.152 $Y=1.487
+ $X2=7.175 $Y2=1.765
r221 31 33 35.5117 $w=2.09e-07 $l=1.54396e-07 $layer=POLY_cond $X=7.152 $Y=1.487
+ $X2=7.115 $Y2=1.35
r222 31 32 61.0776 $w=2.75e-07 $l=2.8e-07 $layer=POLY_cond $X=7.04 $Y=1.487
+ $X2=6.76 $Y2=1.487
r223 28 87 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.685 $Y=1.35
+ $X2=6.685 $Y2=1.557
r224 28 30 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.685 $Y=1.35
+ $X2=6.685 $Y2=0.865
r225 25 86 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.67 $Y=1.765
+ $X2=6.67 $Y2=1.557
r226 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.67 $Y=1.765
+ $X2=6.67 $Y2=2.4
r227 22 84 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.22 $Y=1.765
+ $X2=6.22 $Y2=1.557
r228 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.22 $Y=1.765
+ $X2=6.22 $Y2=2.4
r229 19 83 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.115 $Y=1.35
+ $X2=6.115 $Y2=1.557
r230 19 21 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.115 $Y=1.35
+ $X2=6.115 $Y2=0.865
r231 16 81 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.695 $Y=1.765
+ $X2=5.695 $Y2=1.557
r232 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.695 $Y=1.765
+ $X2=5.695 $Y2=2.4
r233 13 80 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.68 $Y=1.35
+ $X2=5.68 $Y2=1.557
r234 13 15 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.68 $Y=1.35
+ $X2=5.68 $Y2=0.865
r235 4 79 300 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=2 $X=4.29
+ $Y=1.935 $X2=4.465 $Y2=2.115
r236 3 77 300 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=2 $X=1.98
+ $Y=1.935 $X2=2.13 $Y2=2.115
r237 2 73 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.935 $X2=0.73 $Y2=2.11
r238 2 46 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.935 $X2=0.73 $Y2=2.79
r239 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.625 $X2=0.71 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 39 41 43 47
+ 49 54 62 67 72 81 84 89 92 96
r96 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r97 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r98 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r99 85 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 84 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r102 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r103 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r104 76 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r105 76 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r106 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r107 73 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.61 $Y=3.33
+ $X2=6.485 $Y2=3.33
r108 73 75 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.61 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 72 95 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=7.497 $Y2=3.33
r110 72 75 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=6.96 $Y2=3.33
r111 71 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r112 71 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r113 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r114 68 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=3.33
+ $X2=5.465 $Y2=3.33
r115 68 70 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.63 $Y=3.33 $X2=6
+ $Y2=3.33
r116 67 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.36 $Y=3.33
+ $X2=6.485 $Y2=3.33
r117 67 70 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.36 $Y=3.33 $X2=6
+ $Y2=3.33
r118 66 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 63 84 13.8148 $w=1.7e-07 $l=3.58e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=3.272 $Y2=3.33
r121 63 65 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 62 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.465 $Y2=3.33
r123 62 65 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.04 $Y2=3.33
r124 61 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r126 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r127 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r130 55 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.22 $Y2=3.33
r131 55 57 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r132 54 84 13.8148 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.272 $Y2=3.33
r133 54 60 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 53 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r135 53 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r136 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r137 50 78 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r138 50 52 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r139 49 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.22 $Y2=3.33
r140 49 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r141 47 66 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=5.04 $Y2=3.33
r142 47 85 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r143 43 46 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=7.44 $Y=2.115
+ $X2=7.44 $Y2=2.815
r144 41 95 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.44 $Y=3.245
+ $X2=7.497 $Y2=3.33
r145 41 46 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.44 $Y=3.245
+ $X2=7.44 $Y2=2.815
r146 37 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=3.245
+ $X2=6.485 $Y2=3.33
r147 37 39 41.027 $w=2.48e-07 $l=8.9e-07 $layer=LI1_cond $X=6.485 $Y=3.245
+ $X2=6.485 $Y2=2.355
r148 33 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=3.245
+ $X2=5.465 $Y2=3.33
r149 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.465 $Y=3.245
+ $X2=5.465 $Y2=2.415
r150 29 84 2.90666 $w=7.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.272 $Y=3.245
+ $X2=3.272 $Y2=3.33
r151 29 31 13.2154 $w=7.13e-07 $l=7.9e-07 $layer=LI1_cond $X=3.272 $Y=3.245
+ $X2=3.272 $Y2=2.455
r152 25 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r153 25 27 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.455
r154 21 24 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.24 $Y=2.115
+ $X2=0.24 $Y2=2.795
r155 19 78 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r156 19 24 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.795
r157 6 46 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.84 $X2=7.4 $Y2=2.815
r158 6 43 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.84 $X2=7.4 $Y2=2.115
r159 5 39 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=6.295
+ $Y=1.84 $X2=6.445 $Y2=2.355
r160 4 35 300 $w=1.7e-07 $l=5.71314e-07 $layer=licon1_PDIFF $count=2 $X=5.265
+ $Y=1.935 $X2=5.465 $Y2=2.415
r161 3 31 150 $w=1.7e-07 $l=8.56402e-07 $layer=licon1_PDIFF $count=4 $X=2.88
+ $Y=1.935 $X2=3.515 $Y2=2.455
r162 2 27 300 $w=1.7e-07 $l=5.90254e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.935 $X2=1.18 $Y2=2.455
r163 1 24 400 $w=1.7e-07 $l=9.29677e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.935 $X2=0.28 $Y2=2.795
r164 1 21 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.935 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%A_297_387# 1 2 9 11 12 15
r26 13 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.58 $Y=2.905
+ $X2=2.58 $Y2=2.415
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=2.99
+ $X2=2.58 $Y2=2.905
r28 11 12 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.415 $Y=2.99
+ $X2=1.845 $Y2=2.99
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.68 $Y=2.905
+ $X2=1.845 $Y2=2.99
r30 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.68 $Y=2.905 $X2=1.68
+ $Y2=2.415
r31 2 15 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=2.43
+ $Y=1.935 $X2=2.58 $Y2=2.415
r32 1 9 300 $w=1.7e-07 $l=5.6921e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.935 $X2=1.68 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%A_763_387# 1 2 9 11 12 15
c20 11 0 1.23775e-19 $X=4.8 $Y=2.99
r21 13 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.965 $Y=2.905
+ $X2=4.965 $Y2=2.415
r22 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.8 $Y=2.99
+ $X2=4.965 $Y2=2.905
r23 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.8 $Y=2.99 $X2=4.13
+ $Y2=2.99
r24 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.965 $Y=2.905
+ $X2=4.13 $Y2=2.99
r25 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=3.965 $Y=2.905
+ $X2=3.965 $Y2=2.415
r26 2 15 300 $w=1.7e-07 $l=5.71314e-07 $layer=licon1_PDIFF $count=2 $X=4.765
+ $Y=1.935 $X2=4.965 $Y2=2.415
r27 1 9 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=3.815
+ $Y=1.935 $X2=3.965 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%X 1 2 3 4 15 17 19 21 22 23 27 33 37 38 40
+ 44
c71 15 0 1.46284e-19 $X=5.9 $Y=0.64
r72 41 43 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=6.95 $Y=1.935 $X2=6.95
+ $Y2=1.985
r73 39 44 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.115 $Y=1.665
+ $X2=7.44 $Y2=1.665
r74 38 41 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=1.665
+ $X2=6.95 $Y2=1.935
r75 38 40 4.31382 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.95 $Y=1.665
+ $X2=6.95 $Y2=1.55
r76 38 39 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.95 $Y=1.665
+ $X2=7.115 $Y2=1.665
r77 31 43 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6.95 $Y=2.02
+ $X2=6.95 $Y2=1.985
r78 31 33 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=6.95 $Y=2.02
+ $X2=6.95 $Y2=2.815
r79 29 37 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.925 $Y=1.18
+ $X2=6.9 $Y2=1.095
r80 29 40 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=6.925 $Y=1.18
+ $X2=6.925 $Y2=1.55
r81 25 37 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.9 $Y=1.01 $X2=6.9
+ $Y2=1.095
r82 25 27 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.9 $Y=1.01 $X2=6.9
+ $Y2=0.64
r83 24 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.16 $Y=1.935
+ $X2=5.995 $Y2=1.935
r84 23 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=1.935
+ $X2=6.95 $Y2=1.935
r85 23 24 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.785 $Y=1.935
+ $X2=6.16 $Y2=1.935
r86 21 37 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.735 $Y=1.095
+ $X2=6.9 $Y2=1.095
r87 21 22 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.735 $Y=1.095
+ $X2=5.985 $Y2=1.095
r88 17 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.995 $Y=2.02
+ $X2=5.995 $Y2=1.935
r89 17 19 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=5.995 $Y=2.02
+ $X2=5.995 $Y2=2.815
r90 13 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.86 $Y=1.01
+ $X2=5.985 $Y2=1.095
r91 13 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=5.86 $Y=1.01
+ $X2=5.86 $Y2=0.64
r92 4 43 400 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.95 $Y2=1.985
r93 4 33 400 $w=1.7e-07 $l=1.07261e-06 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.95 $Y2=2.815
r94 3 36 400 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=5.77 $Y=1.84
+ $X2=5.995 $Y2=2.015
r95 3 19 400 $w=1.7e-07 $l=1.08167e-06 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.84 $X2=5.995 $Y2=2.815
r96 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.76
+ $Y=0.495 $X2=6.9 $Y2=0.64
r97 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.755
+ $Y=0.495 $X2=5.9 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%A_27_125# 1 2 3 4 15 17 18 21 23 27 29 33 35
+ 36
c68 29 0 1.98018e-19 $X=2.84 $Y=0.37
r69 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.005 $Y=0.455
+ $X2=3.005 $Y2=0.77
r70 30 36 8.61065 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=2.305 $Y=0.37
+ $X2=2.14 $Y2=0.36
r71 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.84 $Y=0.37
+ $X2=3.005 $Y2=0.455
r72 29 30 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.84 $Y=0.37
+ $X2=2.305 $Y2=0.37
r73 25 36 0.89609 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.14 $Y=0.455
+ $X2=2.14 $Y2=0.36
r74 25 27 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.14 $Y=0.455
+ $X2=2.14 $Y2=0.77
r75 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0.35
+ $X2=1.14 $Y2=0.35
r76 23 36 8.61065 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=1.975 $Y=0.35
+ $X2=2.14 $Y2=0.36
r77 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=0.35
+ $X2=1.305 $Y2=0.35
r78 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.435
+ $X2=1.14 $Y2=0.35
r79 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.14 $Y=0.435
+ $X2=1.14 $Y2=0.77
r80 17 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0.35
+ $X2=1.14 $Y2=0.35
r81 17 18 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.975 $Y=0.35
+ $X2=0.365 $Y2=0.35
r82 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.435
+ $X2=0.365 $Y2=0.35
r83 13 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=0.435
+ $X2=0.24 $Y2=0.77
r84 4 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.625 $X2=3.005 $Y2=0.77
r85 3 27 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.625 $X2=2.14 $Y2=0.77
r86 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.625 $X2=1.14 $Y2=0.77
r87 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.625 $X2=0.28 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%A_300_125# 1 2 3 4 13 15 17 21 23 27 29 31
+ 33 38 39
c69 33 0 3.38411e-20 $X=4.89 $Y=0.755
c70 27 0 1.38543e-19 $X=4.025 $Y=0.75
c71 15 0 1.70191e-19 $X=1.64 $Y=0.77
r72 31 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.01 $X2=4.93
+ $Y2=1.095
r73 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.93 $Y=1.01
+ $X2=4.93 $Y2=0.755
r74 30 39 5.29182 $w=1.7e-07 $l=1.08995e-07 $layer=LI1_cond $X=4.115 $Y=1.095
+ $X2=4.027 $Y2=1.142
r75 29 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.805 $Y=1.095
+ $X2=4.93 $Y2=1.095
r76 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.805 $Y=1.095
+ $X2=4.115 $Y2=1.095
r77 25 39 1.23839 $w=1.75e-07 $l=1.32e-07 $layer=LI1_cond $X=4.027 $Y=1.01
+ $X2=4.027 $Y2=1.142
r78 25 27 16.4779 $w=1.73e-07 $l=2.6e-07 $layer=LI1_cond $X=4.027 $Y=1.01
+ $X2=4.027 $Y2=0.75
r79 24 38 4.85493 $w=2.1e-07 $l=1.51687e-07 $layer=LI1_cond $X=2.74 $Y=1.19
+ $X2=2.607 $Y2=1.15
r80 23 39 5.29182 $w=1.7e-07 $l=1.08374e-07 $layer=LI1_cond $X=3.94 $Y=1.19
+ $X2=4.027 $Y2=1.142
r81 23 24 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=3.94 $Y=1.19
+ $X2=2.74 $Y2=1.19
r82 19 38 1.61074 $w=1.95e-07 $l=1.41421e-07 $layer=LI1_cond $X=2.572 $Y=1.025
+ $X2=2.607 $Y2=1.15
r83 19 21 12.7972 $w=1.93e-07 $l=2.25e-07 $layer=LI1_cond $X=2.572 $Y=1.025
+ $X2=2.572 $Y2=0.8
r84 18 36 3.95903 $w=2.5e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.805 $Y=1.15
+ $X2=1.64 $Y2=1.155
r85 17 38 4.85493 $w=2.1e-07 $l=1.32e-07 $layer=LI1_cond $X=2.475 $Y=1.15
+ $X2=2.607 $Y2=1.15
r86 17 18 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=1.15
+ $X2=1.805 $Y2=1.15
r87 13 36 3.0275 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=1.64 $Y=1.025 $X2=1.64
+ $Y2=1.155
r88 13 15 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.64 $Y=1.025
+ $X2=1.64 $Y2=0.77
r89 4 41 182 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_NDIFF $count=1 $X=4.75
+ $Y=0.595 $X2=4.89 $Y2=1.095
r90 4 33 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.75
+ $Y=0.595 $X2=4.89 $Y2=0.755
r91 3 27 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.595 $X2=4.025 $Y2=0.75
r92 2 38 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.625 $X2=2.57 $Y2=1.14
r93 2 21 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.625 $X2=2.57 $Y2=0.8
r94 1 36 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.625 $X2=1.64 $Y2=1.12
r95 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.625 $X2=1.64 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_4%VGND 1 2 3 4 5 18 22 26 32 34 36 39 40 42 43
+ 44 46 61 65 71 74 78
r91 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r92 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r93 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r94 69 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r95 69 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r96 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r97 66 74 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.565 $Y=0 $X2=6.365
+ $Y2=0
r98 66 68 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.565 $Y=0 $X2=6.96
+ $Y2=0
r99 65 77 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.235 $Y=0 $X2=7.457
+ $Y2=0
r100 65 68 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.235 $Y=0
+ $X2=6.96 $Y2=0
r101 64 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r102 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r103 61 74 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.165 $Y=0 $X2=6.365
+ $Y2=0
r104 61 63 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=0 $X2=6
+ $Y2=0
r105 60 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r106 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r107 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r108 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r109 54 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.595
+ $Y2=0
r110 54 56 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=4.08
+ $Y2=0
r111 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r112 52 53 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r113 49 53 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=3.12 $Y2=0
r114 48 52 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.12
+ $Y2=0
r115 48 49 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r116 46 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.595
+ $Y2=0
r117 46 52 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.12
+ $Y2=0
r118 44 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r119 44 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r120 42 59 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.235 $Y=0
+ $X2=5.04 $Y2=0
r121 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.4
+ $Y2=0
r122 41 63 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=6
+ $Y2=0
r123 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.4
+ $Y2=0
r124 39 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=4.08 $Y2=0
r125 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=0 $X2=4.46
+ $Y2=0
r126 38 59 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.625 $Y=0
+ $X2=5.04 $Y2=0
r127 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.46
+ $Y2=0
r128 34 77 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.4 $Y=0.085
+ $X2=7.457 $Y2=0
r129 34 36 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=7.4 $Y=0.085
+ $X2=7.4 $Y2=0.64
r130 30 74 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.365 $Y=0.085
+ $X2=6.365 $Y2=0
r131 30 32 15.9901 $w=3.98e-07 $l=5.55e-07 $layer=LI1_cond $X=6.365 $Y=0.085
+ $X2=6.365 $Y2=0.64
r132 26 28 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=5.4 $Y=0.64
+ $X2=5.4 $Y2=1.055
r133 24 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=0.085 $X2=5.4
+ $Y2=0
r134 24 26 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=5.4 $Y=0.085
+ $X2=5.4 $Y2=0.64
r135 20 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0
r136 20 22 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0.745
r137 16 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=0.085
+ $X2=3.595 $Y2=0
r138 16 18 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=3.595 $Y=0.085
+ $X2=3.595 $Y2=0.755
r139 5 36 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.19
+ $Y=0.495 $X2=7.4 $Y2=0.64
r140 4 32 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=6.19
+ $Y=0.495 $X2=6.365 $Y2=0.64
r141 3 28 182 $w=1.7e-07 $l=5.59285e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.595 $X2=5.4 $Y2=1.055
r142 3 26 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.595 $X2=5.4 $Y2=0.64
r143 2 22 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.32
+ $Y=0.595 $X2=4.46 $Y2=0.745
r144 1 18 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.595 $X2=3.595 $Y2=0.755
.ends

