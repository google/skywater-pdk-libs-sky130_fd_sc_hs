* File: sky130_fd_sc_hs__ha_1.pex.spice
* Created: Tue Sep  1 20:06:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__HA_1%A_83_260# 1 2 9 11 13 14 15 16 18 19 25 29
c59 25 0 5.39611e-20 $X=1.235 $Y=1.105
c60 16 0 3.29783e-20 $X=1.07 $Y=1.215
c61 2 0 1.20626e-19 $X=1.425 $Y=1.96
r62 29 32 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.575 $Y=2.395
+ $X2=1.575 $Y2=2.555
r63 25 27 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.235 $Y=1.105
+ $X2=1.235 $Y2=1.215
r64 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.465 $X2=0.69 $Y2=1.465
r65 20 22 11.0909 $w=2.75e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=1.215
+ $X2=0.69 $Y2=1.465
r66 18 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=2.395
+ $X2=1.575 $Y2=2.395
r67 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.41 $Y=2.395
+ $X2=0.855 $Y2=2.395
r68 17 20 3.55113 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=1.215
+ $X2=0.69 $Y2=1.215
r69 16 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=1.215
+ $X2=1.235 $Y2=1.215
r70 16 17 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.07 $Y=1.215
+ $X2=0.855 $Y2=1.215
r71 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.77 $Y=2.31
+ $X2=0.855 $Y2=2.395
r72 14 22 9.08745 $w=2.75e-07 $l=2.0106e-07 $layer=LI1_cond $X=0.77 $Y=1.63
+ $X2=0.69 $Y2=1.465
r73 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.77 $Y=1.63
+ $X2=0.77 $Y2=2.31
r74 11 23 56.8427 $w=3.64e-07 $l=3.59166e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.635 $Y2=1.465
r75 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r76 7 23 38.9663 $w=3.64e-07 $l=2.24332e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.635 $Y2=1.465
r77 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
r78 2 32 600 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.96 $X2=1.575 $Y2=2.555
r79 1 25 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.93 $X2=1.235 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_HS__HA_1%A_239_294# 1 2 7 9 12 14 16 17 19 22 25 26 29
+ 33 36 37 39 44
c112 37 0 1.20589e-19 $X=3.64 $Y=1.515
c113 29 0 9.69512e-20 $X=3.185 $Y=0.74
c114 22 0 2.42375e-19 $X=1.36 $Y=1.635
c115 12 0 1.11764e-19 $X=1.45 $Y=0.97
r116 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.515 $X2=4.21 $Y2=1.515
r117 37 43 3.39238 $w=3.3e-07 $l=2.995e-07 $layer=LI1_cond $X=3.64 $Y=1.515
+ $X2=3.555 $Y2=1.255
r118 37 39 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=3.64 $Y=1.515
+ $X2=4.21 $Y2=1.515
r119 36 44 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=3.555 $Y=1.97
+ $X2=3.5 $Y2=2.055
r120 35 43 3.78059 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=3.555 $Y=1.68
+ $X2=3.555 $Y2=1.255
r121 35 36 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.555 $Y=1.68
+ $X2=3.555 $Y2=1.97
r122 31 44 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=2.14 $X2=3.5
+ $Y2=2.055
r123 31 33 5.14483 $w=2.78e-07 $l=1.25e-07 $layer=LI1_cond $X=3.5 $Y=2.14
+ $X2=3.5 $Y2=2.265
r124 27 43 15.7832 $w=2.86e-07 $l=3.7e-07 $layer=LI1_cond $X=3.185 $Y=1.255
+ $X2=3.555 $Y2=1.255
r125 27 29 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.185 $Y=1.085
+ $X2=3.185 $Y2=0.74
r126 25 44 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.36 $Y=2.055
+ $X2=3.5 $Y2=2.055
r127 25 26 119.717 $w=1.68e-07 $l=1.835e-06 $layer=LI1_cond $X=3.36 $Y=2.055
+ $X2=1.525 $Y2=2.055
r128 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.36
+ $Y=1.635 $X2=1.36 $Y2=1.635
r129 20 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.36 $Y=1.97
+ $X2=1.525 $Y2=2.055
r130 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.36 $Y=1.97
+ $X2=1.36 $Y2=1.635
r131 17 40 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=4.26 $Y=1.35
+ $X2=4.21 $Y2=1.515
r132 17 19 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.26 $Y=1.35
+ $X2=4.26 $Y2=0.865
r133 14 40 52.2586 $w=2.99e-07 $l=2.69258e-07 $layer=POLY_cond $X=4.25 $Y=1.765
+ $X2=4.21 $Y2=1.515
r134 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.25 $Y=1.765
+ $X2=4.25 $Y2=2.4
r135 10 23 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.45 $Y=1.47
+ $X2=1.36 $Y2=1.635
r136 10 12 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.45 $Y=1.47 $X2=1.45
+ $Y2=0.97
r137 7 23 52.2586 $w=2.99e-07 $l=2.54951e-07 $layer=POLY_cond $X=1.35 $Y=1.885
+ $X2=1.36 $Y2=1.635
r138 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.35 $Y=1.885
+ $X2=1.35 $Y2=2.38
r139 2 33 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.325
+ $Y=2.12 $X2=3.475 $Y2=2.265
r140 1 29 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.04
+ $Y=0.595 $X2=3.185 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__HA_1%B 1 3 6 9 10 12 15 23 24 30 33
c65 24 0 1.87829e-19 $X=3.12 $Y=1.665
c66 23 0 1.35157e-19 $X=2.095 $Y=1.635
c67 6 0 2.89045e-19 $X=1.88 $Y=0.97
r68 28 30 19.726 $w=2.81e-07 $l=1.15e-07 $layer=POLY_cond $X=3.135 $Y=1.635
+ $X2=3.25 $Y2=1.635
r69 24 33 5.94304 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.12 $Y=1.635
+ $X2=2.97 $Y2=1.635
r70 24 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.135
+ $Y=1.635 $X2=3.135 $Y2=1.635
r71 23 33 40.3355 $w=2.48e-07 $l=8.75e-07 $layer=LI1_cond $X=2.095 $Y=1.675
+ $X2=2.97 $Y2=1.675
r72 20 23 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=1.635
+ $X2=2.095 $Y2=1.635
r73 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.635 $X2=1.93 $Y2=1.635
r74 13 30 25.7295 $w=2.81e-07 $l=2.2798e-07 $layer=POLY_cond $X=3.4 $Y=1.47
+ $X2=3.25 $Y2=1.635
r75 13 15 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.4 $Y=1.47 $X2=3.4
+ $Y2=0.915
r76 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.25 $Y=2.045
+ $X2=3.25 $Y2=2.54
r77 9 10 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.25 $Y=1.955 $X2=3.25
+ $Y2=2.045
r78 8 30 13.2092 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.8 $X2=3.25
+ $Y2=1.635
r79 8 9 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=3.25 $Y=1.8 $X2=3.25
+ $Y2=1.955
r80 4 21 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=1.88 $Y=1.47
+ $X2=1.93 $Y2=1.635
r81 4 6 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.88 $Y=1.47 $X2=1.88
+ $Y2=0.97
r82 1 21 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.855 $Y=1.885
+ $X2=1.93 $Y2=1.635
r83 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.855 $Y=1.885
+ $X2=1.855 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__HA_1%A 4 5 6 7 9 10 12 14 16 18 20 22 26
c72 26 0 9.52888e-20 $X=2.615 $Y=0.42
c73 22 0 9.69512e-20 $X=2.557 $Y=0.18
c74 18 0 1.87829e-19 $X=3.76 $Y=0.915
c75 16 0 1.11259e-19 $X=3.76 $Y=1.86
r76 25 27 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=2.557 $Y=0.42
+ $X2=2.557 $Y2=0.585
r77 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=0.42 $X2=2.615 $Y2=0.42
r78 22 25 29.9948 $w=4.45e-07 $l=2.4e-07 $layer=POLY_cond $X=2.557 $Y=0.18
+ $X2=2.557 $Y2=0.42
r79 20 26 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.615 $Y=0.555
+ $X2=2.615 $Y2=0.42
r80 16 18 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=3.76 $Y=1.86
+ $X2=3.76 $Y2=0.915
r81 15 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.76 $Y=0.255
+ $X2=3.76 $Y2=0.915
r82 12 16 41.2824 $w=2.16e-07 $l=2.12897e-07 $layer=POLY_cond $X=3.7 $Y=2.045
+ $X2=3.76 $Y2=1.86
r83 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.7 $Y=2.045 $X2=3.7
+ $Y2=2.54
r84 11 22 28.4889 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.78 $Y=0.18
+ $X2=2.557 $Y2=0.18
r85 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.685 $Y=0.18
+ $X2=3.76 $Y2=0.255
r86 10 11 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=3.685 $Y=0.18
+ $X2=2.78 $Y2=0.18
r87 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.885
+ $X2=2.425 $Y2=2.46
r88 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.425 $Y=1.795 $X2=2.425
+ $Y2=1.885
r89 5 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.425 $Y=1.5 $X2=2.425
+ $Y2=1.41
r90 5 6 114.669 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=2.425 $Y=1.5
+ $X2=2.425 $Y2=1.795
r91 4 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.41 $Y=1.015
+ $X2=2.41 $Y2=1.41
r92 4 27 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.41 $Y=1.015
+ $X2=2.41 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HS__HA_1%SUM 1 2 7 8 9 10 11 12 13 30 40
r22 23 30 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=0.28 $Y=0.965 $X2=0.28
+ $Y2=0.925
r23 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=2.405
+ $X2=0.28 $Y2=2.775
r24 11 40 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=0.28 $Y=1.967
+ $X2=0.28 $Y2=1.985
r25 11 51 6.01134 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=0.28 $Y=1.967
+ $X2=0.28 $Y2=1.82
r26 11 12 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=0.28 $Y=2.052
+ $X2=0.28 $Y2=2.405
r27 11 40 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=0.28 $Y=2.052
+ $X2=0.28 $Y2=1.985
r28 10 51 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=0.235 $Y=1.665
+ $X2=0.235 $Y2=1.82
r29 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r30 9 49 7.92305 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.13
r31 8 49 5.87165 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=0.28 $Y=0.987
+ $X2=0.28 $Y2=1.13
r32 8 23 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=0.28 $Y=0.987
+ $X2=0.28 $Y2=0.965
r33 8 30 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=0.28 $Y=0.902
+ $X2=0.28 $Y2=0.925
r34 7 8 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=0.28 $Y=0.515 $X2=0.28
+ $Y2=0.902
r35 2 13 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r36 2 40 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r37 1 7 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__HA_1%VPWR 1 2 3 12 16 20 23 24 25 27 32 42 43 46 51
c61 1 0 1.21749e-19 $X=0.58 $Y=1.84
r62 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 47 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 46 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r67 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r68 40 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r70 37 51 13.7128 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=3.19 $Y=3.33
+ $X2=2.837 $Y2=3.33
r71 37 39 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.19 $Y=3.33 $X2=3.6
+ $Y2=3.33
r72 36 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 33 46 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=0.91 $Y2=3.33
r75 33 35 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 32 51 13.7128 $w=1.7e-07 $l=3.52e-07 $layer=LI1_cond $X=2.485 $Y=3.33
+ $X2=2.837 $Y2=3.33
r77 32 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 30 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 27 46 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.91 $Y2=3.33
r81 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r82 25 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r83 25 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 23 39 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=3.33 $X2=3.6
+ $Y2=3.33
r85 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=3.33
+ $X2=3.975 $Y2=3.33
r86 22 42 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.14 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=3.33
+ $X2=3.975 $Y2=3.33
r88 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=3.245
+ $X2=3.975 $Y2=3.33
r89 18 20 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=3.975 $Y=3.245
+ $X2=3.975 $Y2=2.265
r90 14 51 2.87722 $w=7.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.837 $Y=3.245
+ $X2=2.837 $Y2=3.33
r91 14 16 14.4208 $w=7.03e-07 $l=8.5e-07 $layer=LI1_cond $X=2.837 $Y=3.245
+ $X2=2.837 $Y2=2.395
r92 10 46 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=3.245
+ $X2=0.91 $Y2=3.33
r93 10 12 9.52808 $w=5.88e-07 $l=4.7e-07 $layer=LI1_cond $X=0.91 $Y=3.245
+ $X2=0.91 $Y2=2.775
r94 3 20 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=3.775
+ $Y=2.12 $X2=3.975 $Y2=2.265
r95 2 16 150 $w=1.7e-07 $l=7.0993e-07 $layer=licon1_PDIFF $count=4 $X=2.5
+ $Y=1.96 $X2=3.025 $Y2=2.395
r96 1 12 600 $w=1.7e-07 $l=1.09184e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.92 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_HS__HA_1%COUT 1 2 9 13 14 15 16 30
c24 14 0 1.11259e-19 $X=4.56 $Y=2.035
r25 15 16 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=4.512 $Y=2.405
+ $X2=4.512 $Y2=2.775
r26 14 21 1.45122 $w=4.03e-07 $l=5.1e-08 $layer=LI1_cond $X=4.512 $Y=2.001
+ $X2=4.512 $Y2=2.052
r27 14 30 8.27043 $w=4.03e-07 $l=1.51e-07 $layer=LI1_cond $X=4.512 $Y=2.001
+ $X2=4.512 $Y2=1.85
r28 14 15 9.07727 $w=4.03e-07 $l=3.19e-07 $layer=LI1_cond $X=4.512 $Y=2.086
+ $X2=4.512 $Y2=2.405
r29 14 21 0.967483 $w=4.03e-07 $l=3.4e-08 $layer=LI1_cond $X=4.512 $Y=2.086
+ $X2=4.512 $Y2=2.052
r30 13 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.63 $Y=1.18
+ $X2=4.63 $Y2=1.85
r31 7 13 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=4.512 $Y=0.978
+ $X2=4.512 $Y2=1.18
r32 7 9 9.61792 $w=4.03e-07 $l=3.38e-07 $layer=LI1_cond $X=4.512 $Y=0.978
+ $X2=4.512 $Y2=0.64
r33 2 14 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.84 $X2=4.475 $Y2=2.015
r34 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.84 $X2=4.475 $Y2=2.815
r35 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.335
+ $Y=0.495 $X2=4.475 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_HS__HA_1%VGND 1 2 3 12 16 20 23 24 25 27 32 45 46 49 52
r55 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r58 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r59 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r60 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r61 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r62 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r63 37 52 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.105
+ $Y2=0
r64 37 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.64
+ $Y2=0
r65 36 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r66 36 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r67 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 33 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.75
+ $Y2=0
r69 33 35 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.68
+ $Y2=0
r70 32 52 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.105
+ $Y2=0
r71 32 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.68
+ $Y2=0
r72 30 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r73 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r74 27 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.75
+ $Y2=0
r75 27 29 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r76 25 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r77 25 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r78 23 42 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.6
+ $Y2=0
r79 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.975
+ $Y2=0
r80 22 45 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.56
+ $Y2=0
r81 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=3.975
+ $Y2=0
r82 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=0.085
+ $X2=3.975 $Y2=0
r83 18 20 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.975 $Y=0.085
+ $X2=3.975 $Y2=0.72
r84 14 52 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r85 14 16 23.3781 $w=3.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.795
r86 10 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r87 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.515
r88 3 20 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.835
+ $Y=0.595 $X2=3.975 $Y2=0.72
r89 2 16 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.65 $X2=2.105 $Y2=0.795
r90 1 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__HA_1%A_305_130# 1 2 9 11 12 14
c28 12 0 7.8786e-20 $X=1.75 $Y=1.215
c29 9 0 1.39795e-19 $X=1.665 $Y=0.795
r30 14 16 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.625 $Y=1.095
+ $X2=2.625 $Y2=1.215
r31 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=1.215
+ $X2=2.625 $Y2=1.215
r32 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.46 $Y=1.215
+ $X2=1.75 $Y2=1.215
r33 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.665 $Y=1.13
+ $X2=1.75 $Y2=1.215
r34 7 9 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=1.13
+ $X2=1.665 $Y2=0.795
r35 2 14 182 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.695 $X2=2.625 $Y2=1.095
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.525
+ $Y=0.65 $X2=1.665 $Y2=0.795
.ends

