* File: sky130_fd_sc_hs__or4b_4.pxi.spice
* Created: Thu Aug 27 21:07:20 2020
* 
x_PM_SKY130_FD_SC_HS__OR4B_4%B N_B_c_130_n N_B_M1020_g N_B_c_140_n N_B_M1006_g
+ N_B_c_131_n N_B_c_142_n N_B_M1011_g N_B_c_132_n N_B_c_133_n N_B_c_134_n B B
+ N_B_c_135_n N_B_c_136_n N_B_c_137_n N_B_c_138_n PM_SKY130_FD_SC_HS__OR4B_4%B
x_PM_SKY130_FD_SC_HS__OR4B_4%A N_A_c_210_n N_A_M1007_g N_A_M1021_g N_A_c_211_n
+ N_A_M1010_g A N_A_c_209_n PM_SKY130_FD_SC_HS__OR4B_4%A
x_PM_SKY130_FD_SC_HS__OR4B_4%C N_C_M1018_g N_C_c_255_n N_C_c_266_n N_C_M1009_g
+ N_C_c_256_n N_C_c_268_n N_C_M1015_g N_C_c_257_n N_C_c_258_n N_C_c_259_n
+ N_C_c_260_n C N_C_c_261_n N_C_c_262_n N_C_c_263_n N_C_c_264_n
+ PM_SKY130_FD_SC_HS__OR4B_4%C
x_PM_SKY130_FD_SC_HS__OR4B_4%A_563_48# N_A_563_48#_M1016_s N_A_563_48#_M1004_s
+ N_A_563_48#_M1019_g N_A_563_48#_c_356_n N_A_563_48#_M1008_g
+ N_A_563_48#_c_357_n N_A_563_48#_M1012_g N_A_563_48#_c_351_n
+ N_A_563_48#_c_352_n N_A_563_48#_c_353_n N_A_563_48#_c_358_n
+ N_A_563_48#_c_354_n N_A_563_48#_c_360_n N_A_563_48#_c_355_n
+ PM_SKY130_FD_SC_HS__OR4B_4%A_563_48#
x_PM_SKY130_FD_SC_HS__OR4B_4%D_N N_D_N_c_444_n N_D_N_M1016_g N_D_N_c_445_n
+ N_D_N_M1004_g D_N PM_SKY130_FD_SC_HS__OR4B_4%D_N
x_PM_SKY130_FD_SC_HS__OR4B_4%A_27_74# N_A_27_74#_M1020_s N_A_27_74#_M1021_d
+ N_A_27_74#_M1019_d N_A_27_74#_M1008_d N_A_27_74#_M1001_g N_A_27_74#_c_496_n
+ N_A_27_74#_M1000_g N_A_27_74#_M1013_g N_A_27_74#_c_497_n N_A_27_74#_M1002_g
+ N_A_27_74#_c_498_n N_A_27_74#_M1003_g N_A_27_74#_M1014_g N_A_27_74#_c_499_n
+ N_A_27_74#_M1005_g N_A_27_74#_M1017_g N_A_27_74#_c_484_n N_A_27_74#_c_485_n
+ N_A_27_74#_c_486_n N_A_27_74#_c_487_n N_A_27_74#_c_488_n N_A_27_74#_c_489_n
+ N_A_27_74#_c_490_n N_A_27_74#_c_491_n N_A_27_74#_c_492_n N_A_27_74#_c_493_n
+ N_A_27_74#_c_581_p N_A_27_74#_c_512_n N_A_27_74#_c_494_n N_A_27_74#_c_534_n
+ N_A_27_74#_c_495_n PM_SKY130_FD_SC_HS__OR4B_4%A_27_74#
x_PM_SKY130_FD_SC_HS__OR4B_4%A_27_392# N_A_27_392#_M1006_s N_A_27_392#_M1011_s
+ N_A_27_392#_M1015_s N_A_27_392#_c_674_n N_A_27_392#_c_675_n
+ N_A_27_392#_c_676_n N_A_27_392#_c_677_n N_A_27_392#_c_702_n
+ N_A_27_392#_c_678_n N_A_27_392#_c_704_n N_A_27_392#_c_679_n
+ N_A_27_392#_c_680_n N_A_27_392#_c_708_n N_A_27_392#_c_681_n
+ PM_SKY130_FD_SC_HS__OR4B_4%A_27_392#
x_PM_SKY130_FD_SC_HS__OR4B_4%A_116_392# N_A_116_392#_M1006_d
+ N_A_116_392#_M1010_s N_A_116_392#_c_751_n N_A_116_392#_c_747_n
+ N_A_116_392#_c_748_n PM_SKY130_FD_SC_HS__OR4B_4%A_116_392#
x_PM_SKY130_FD_SC_HS__OR4B_4%VPWR N_VPWR_M1007_d N_VPWR_M1004_d N_VPWR_M1002_s
+ N_VPWR_M1005_s N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n N_VPWR_c_774_n
+ N_VPWR_c_775_n VPWR N_VPWR_c_776_n N_VPWR_c_777_n N_VPWR_c_778_n
+ N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n N_VPWR_c_770_n
+ PM_SKY130_FD_SC_HS__OR4B_4%VPWR
x_PM_SKY130_FD_SC_HS__OR4B_4%A_496_392# N_A_496_392#_M1009_d
+ N_A_496_392#_M1012_s N_A_496_392#_c_860_n
+ PM_SKY130_FD_SC_HS__OR4B_4%A_496_392#
x_PM_SKY130_FD_SC_HS__OR4B_4%X N_X_M1001_s N_X_M1014_s N_X_M1000_d N_X_M1003_d
+ N_X_c_873_n N_X_c_880_n N_X_c_881_n N_X_c_874_n N_X_c_875_n N_X_c_882_n
+ N_X_c_876_n N_X_c_883_n N_X_c_884_n N_X_c_877_n N_X_c_878_n N_X_c_879_n X X
+ PM_SKY130_FD_SC_HS__OR4B_4%X
x_PM_SKY130_FD_SC_HS__OR4B_4%VGND N_VGND_M1020_d N_VGND_M1018_d N_VGND_M1016_d
+ N_VGND_M1013_d N_VGND_M1017_d N_VGND_c_950_n N_VGND_c_951_n N_VGND_c_952_n
+ N_VGND_c_953_n N_VGND_c_954_n N_VGND_c_955_n VGND N_VGND_c_956_n
+ N_VGND_c_957_n N_VGND_c_958_n N_VGND_c_959_n N_VGND_c_960_n N_VGND_c_961_n
+ N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n N_VGND_c_965_n
+ PM_SKY130_FD_SC_HS__OR4B_4%VGND
cc_1 VNB N_B_c_130_n 0.0093615f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.795
cc_2 VNB N_B_c_131_n 0.00657435f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.795
cc_3 VNB N_B_c_132_n 0.0160839f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=1.195
cc_4 VNB N_B_c_133_n 0.00321396f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.195
cc_5 VNB N_B_c_134_n 0.0385296f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.385
cc_6 VNB N_B_c_135_n 0.0356219f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.385
cc_7 VNB N_B_c_136_n 0.0226215f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.22
cc_8 VNB N_B_c_137_n 0.023141f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.33
cc_9 VNB N_B_c_138_n 0.00809179f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.33
cc_10 VNB N_A_M1021_g 0.0372567f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_11 VNB A 0.00179937f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.885
cc_12 VNB N_A_c_209_n 0.0350539f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.195
cc_13 VNB N_C_c_255_n 0.00533349f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_14 VNB N_C_c_256_n 0.011669f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.795
cc_15 VNB N_C_c_257_n 0.00936312f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=1.195
cc_16 VNB N_C_c_258_n 0.00512252f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.195
cc_17 VNB N_C_c_259_n 0.00419907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C_c_260_n 0.00451087f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.385
cc_19 VNB N_C_c_261_n 0.0281686f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_C_c_262_n 0.0217009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_c_263_n 0.0492861f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.55
cc_22 VNB N_C_c_264_n 0.00824303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_563_48#_M1019_g 0.0330273f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.55
cc_24 VNB N_A_563_48#_c_351_n 0.0528013f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.385
cc_25 VNB N_A_563_48#_c_352_n 0.0505231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_563_48#_c_353_n 0.0128142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_563_48#_c_354_n 0.00345786f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.385
cc_28 VNB N_A_563_48#_c_355_n 0.0253522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_D_N_c_444_n 0.019771f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_30 VNB N_D_N_c_445_n 0.0492085f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_31 VNB D_N 0.00753989f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_32 VNB N_A_27_74#_M1001_g 0.0241971f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.195
cc_33 VNB N_A_27_74#_M1013_g 0.0236719f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_A_27_74#_M1014_g 0.0219571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_M1017_g 0.0292173f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.33
cc_36 VNB N_A_27_74#_c_484_n 0.0185887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_485_n 0.00750337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_486_n 0.00457144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_487_n 0.00237713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_488_n 0.00322465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_489_n 0.00566983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_490_n 0.00384103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_491_n 0.0229281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_74#_c_492_n 0.00151598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_74#_c_493_n 0.00404584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_74#_c_494_n 0.00283535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_495_n 0.1202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VPWR_c_770_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_X_c_873_n 0.00326562f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.195
cc_50 VNB N_X_c_874_n 0.0033499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_X_c_875_n 0.00280894f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_52 VNB N_X_c_876_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.385
cc_53 VNB N_X_c_877_n 3.46234e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.33
cc_54 VNB N_X_c_878_n 0.00140937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_X_c_879_n 0.00224001f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.33
cc_56 VNB N_VGND_c_950_n 0.0097033f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.385
cc_57 VNB N_VGND_c_951_n 0.0067114f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_58 VNB N_VGND_c_952_n 0.00940833f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.385
cc_59 VNB N_VGND_c_953_n 0.00503037f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.55
cc_60 VNB N_VGND_c_954_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_955_n 0.0503969f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.33
cc_62 VNB N_VGND_c_956_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.33
cc_63 VNB N_VGND_c_957_n 0.0366654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_958_n 0.0549039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_959_n 0.0183788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_960_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_961_n 0.00632182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_962_n 0.00661316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_963_n 0.00617178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_964_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_965_n 0.392526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VPB N_B_c_130_n 0.0115096f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.795
cc_73 VPB N_B_c_140_n 0.0295146f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_74 VPB N_B_c_131_n 0.00808706f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.795
cc_75 VPB N_B_c_142_n 0.0230404f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.885
cc_76 VPB N_A_c_210_n 0.0152861f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.55
cc_77 VPB N_A_c_211_n 0.0156703f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_78 VPB A 0.00250427f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.885
cc_79 VPB N_A_c_209_n 0.0338722f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.195
cc_80 VPB N_C_c_255_n 0.0067307f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_81 VPB N_C_c_266_n 0.0232421f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_82 VPB N_C_c_256_n 0.00929514f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.795
cc_83 VPB N_C_c_268_n 0.0260827f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.885
cc_84 VPB N_C_c_264_n 0.00650907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_563_48#_c_356_n 0.0158419f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.885
cc_86 VPB N_A_563_48#_c_357_n 0.0157679f $X=-0.19 $Y=1.66 $X2=1.705 $Y2=1.195
cc_87 VPB N_A_563_48#_c_358_n 0.0277449f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.385
cc_88 VPB N_A_563_48#_c_354_n 0.00437779f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.385
cc_89 VPB N_A_563_48#_c_360_n 0.0130255f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.55
cc_90 VPB N_A_563_48#_c_355_n 0.0343514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_D_N_c_445_n 0.0275893f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_92 VPB N_A_27_74#_c_496_n 0.0163765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_74#_c_497_n 0.0148844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_27_74#_c_498_n 0.0148641f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.385
cc_95 VPB N_A_27_74#_c_499_n 0.018379f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.33
cc_96 VPB N_A_27_74#_c_490_n 0.00139272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_74#_c_495_n 0.0291006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_27_392#_c_674_n 0.0112901f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.795
cc_99 VPB N_A_27_392#_c_675_n 0.035396f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=2.46
cc_100 VPB N_A_27_392#_c_676_n 0.0107646f $X=-0.19 $Y=1.66 $X2=1.705 $Y2=1.195
cc_101 VPB N_A_27_392#_c_677_n 0.00934903f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.195
cc_102 VPB N_A_27_392#_c_678_n 0.00289722f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.385
cc_103 VPB N_A_27_392#_c_679_n 0.0027871f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.385
cc_104 VPB N_A_27_392#_c_680_n 0.00730784f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.55
cc_105 VPB N_A_27_392#_c_681_n 0.00153232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_116_392#_c_747_n 0.00180959f $X=-0.19 $Y=1.66 $X2=1.705 $Y2=1.195
cc_107 VPB N_A_116_392#_c_748_n 0.00289794f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.195
cc_108 VPB N_VPWR_c_771_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.195
cc_109 VPB N_VPWR_c_772_n 0.0157217f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.385
cc_110 VPB N_VPWR_c_773_n 0.00271781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_774_n 0.0118511f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.385
cc_112 VPB N_VPWR_c_775_n 0.0345059f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.22
cc_113 VPB N_VPWR_c_776_n 0.0304099f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.55
cc_114 VPB N_VPWR_c_777_n 0.096139f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.33
cc_115 VPB N_VPWR_c_778_n 0.0182909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_779_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_780_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_781_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_782_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_770_n 0.100608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_496_392#_c_860_n 0.00792862f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.885
cc_122 VPB N_X_c_880_n 0.0016237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_X_c_881_n 0.00243101f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.385
cc_124 VPB N_X_c_882_n 0.00228088f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_125 VPB N_X_c_883_n 0.00233217f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.55
cc_126 VPB N_X_c_884_n 0.00153448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB X 0.0244193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 N_B_c_140_n N_A_c_210_n 0.0213251f $X=0.505 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_129 N_B_c_132_n N_A_M1021_g 0.0129521f $X=1.705 $Y=1.195 $X2=0 $Y2=0
cc_130 N_B_c_133_n N_A_M1021_g 0.00113261f $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_131 N_B_c_134_n N_A_M1021_g 0.00486674f $X=1.87 $Y=1.385 $X2=0 $Y2=0
cc_132 N_B_c_135_n N_A_M1021_g 0.00594475f $X=0.43 $Y=1.385 $X2=0 $Y2=0
cc_133 N_B_c_136_n N_A_M1021_g 0.0243288f $X=0.43 $Y=1.22 $X2=0 $Y2=0
cc_134 N_B_c_138_n N_A_M1021_g 0.00495309f $X=0.835 $Y=1.33 $X2=0 $Y2=0
cc_135 N_B_c_142_n N_A_c_211_n 0.0277294f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_136 N_B_c_131_n A 0.00105466f $X=1.905 $Y=1.795 $X2=0 $Y2=0
cc_137 N_B_c_132_n A 0.0242717f $X=1.705 $Y=1.195 $X2=0 $Y2=0
cc_138 N_B_c_133_n A 0.0040169f $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_139 N_B_c_134_n A 2.74307e-19 $X=1.87 $Y=1.385 $X2=0 $Y2=0
cc_140 N_B_c_135_n A 0.00118781f $X=0.43 $Y=1.385 $X2=0 $Y2=0
cc_141 N_B_c_138_n A 0.00837769f $X=0.835 $Y=1.33 $X2=0 $Y2=0
cc_142 N_B_c_131_n N_A_c_209_n 0.0154069f $X=1.905 $Y=1.795 $X2=0 $Y2=0
cc_143 N_B_c_132_n N_A_c_209_n 0.0102355f $X=1.705 $Y=1.195 $X2=0 $Y2=0
cc_144 N_B_c_133_n N_A_c_209_n 4.35205e-19 $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_145 N_B_c_134_n N_A_c_209_n 0.00658941f $X=1.87 $Y=1.385 $X2=0 $Y2=0
cc_146 N_B_c_135_n N_A_c_209_n 0.0228067f $X=0.43 $Y=1.385 $X2=0 $Y2=0
cc_147 N_B_c_138_n N_A_c_209_n 9.92831e-19 $X=0.835 $Y=1.33 $X2=0 $Y2=0
cc_148 N_B_c_131_n N_C_c_255_n 0.00641167f $X=1.905 $Y=1.795 $X2=0 $Y2=0
cc_149 N_B_c_142_n N_C_c_266_n 0.0277771f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_150 N_B_c_133_n N_C_c_258_n 9.75844e-19 $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_151 N_B_c_133_n N_C_c_261_n 4.1682e-19 $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_152 N_B_c_134_n N_C_c_261_n 0.020758f $X=1.87 $Y=1.385 $X2=0 $Y2=0
cc_153 N_B_c_133_n N_C_c_262_n 0.00280031f $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_154 N_B_c_131_n N_C_c_264_n 0.00540384f $X=1.905 $Y=1.795 $X2=0 $Y2=0
cc_155 N_B_c_133_n N_C_c_264_n 0.023338f $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_156 N_B_c_134_n N_C_c_264_n 0.00114908f $X=1.87 $Y=1.385 $X2=0 $Y2=0
cc_157 N_B_c_133_n N_A_27_74#_M1021_d 0.00359065f $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_158 N_B_c_136_n N_A_27_74#_c_484_n 0.00663104f $X=0.43 $Y=1.22 $X2=0 $Y2=0
cc_159 N_B_c_135_n N_A_27_74#_c_485_n 7.83044e-19 $X=0.43 $Y=1.385 $X2=0 $Y2=0
cc_160 N_B_c_136_n N_A_27_74#_c_485_n 7.15561e-19 $X=0.43 $Y=1.22 $X2=0 $Y2=0
cc_161 N_B_c_137_n N_A_27_74#_c_485_n 0.0253334f $X=0.615 $Y=1.33 $X2=0 $Y2=0
cc_162 N_B_c_132_n N_A_27_74#_c_486_n 0.0304032f $X=1.705 $Y=1.195 $X2=0 $Y2=0
cc_163 N_B_c_133_n N_A_27_74#_c_486_n 0.028164f $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_164 N_B_c_134_n N_A_27_74#_c_486_n 0.00192194f $X=1.87 $Y=1.385 $X2=0 $Y2=0
cc_165 N_B_c_136_n N_A_27_74#_c_487_n 5.79051e-19 $X=0.43 $Y=1.22 $X2=0 $Y2=0
cc_166 N_B_c_138_n N_A_27_74#_c_487_n 0.0304032f $X=0.835 $Y=1.33 $X2=0 $Y2=0
cc_167 N_B_c_136_n N_A_27_74#_c_512_n 0.008978f $X=0.43 $Y=1.22 $X2=0 $Y2=0
cc_168 N_B_c_137_n N_A_27_74#_c_512_n 0.0304032f $X=0.615 $Y=1.33 $X2=0 $Y2=0
cc_169 N_B_c_140_n N_A_27_392#_c_674_n 0.00166528f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_170 N_B_c_135_n N_A_27_392#_c_674_n 0.00304873f $X=0.43 $Y=1.385 $X2=0 $Y2=0
cc_171 N_B_c_137_n N_A_27_392#_c_674_n 0.0153775f $X=0.615 $Y=1.33 $X2=0 $Y2=0
cc_172 N_B_c_140_n N_A_27_392#_c_675_n 0.0105177f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_173 N_B_c_140_n N_A_27_392#_c_676_n 0.0135407f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_174 N_B_c_142_n N_A_27_392#_c_676_n 0.0174766f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_175 N_B_c_132_n N_A_27_392#_c_676_n 0.014507f $X=1.705 $Y=1.195 $X2=0 $Y2=0
cc_176 N_B_c_133_n N_A_27_392#_c_676_n 0.0119479f $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_177 N_B_c_134_n N_A_27_392#_c_676_n 7.48688e-19 $X=1.87 $Y=1.385 $X2=0 $Y2=0
cc_178 N_B_c_137_n N_A_27_392#_c_676_n 0.0163004f $X=0.615 $Y=1.33 $X2=0 $Y2=0
cc_179 N_B_c_133_n N_A_27_392#_c_677_n 8.65747e-19 $X=1.87 $Y=1.195 $X2=0 $Y2=0
cc_180 N_B_c_142_n N_A_27_392#_c_678_n 0.00245875f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_181 N_B_c_140_n N_A_116_392#_c_747_n 0.00172473f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_B_c_142_n N_A_116_392#_c_748_n 0.00712193f $X=1.905 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_B_c_140_n N_VPWR_c_771_n 6.41695e-19 $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_184 N_B_c_142_n N_VPWR_c_771_n 6.11631e-19 $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_185 N_B_c_140_n N_VPWR_c_776_n 0.00445602f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_186 N_B_c_142_n N_VPWR_c_777_n 0.00445602f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_187 N_B_c_140_n N_VPWR_c_770_n 0.00861929f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_188 N_B_c_142_n N_VPWR_c_770_n 0.0085938f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_189 N_B_c_136_n N_VGND_c_950_n 0.0047684f $X=0.43 $Y=1.22 $X2=0 $Y2=0
cc_190 N_B_c_136_n N_VGND_c_956_n 0.00434272f $X=0.43 $Y=1.22 $X2=0 $Y2=0
cc_191 N_B_c_136_n N_VGND_c_965_n 0.00435167f $X=0.43 $Y=1.22 $X2=0 $Y2=0
cc_192 N_A_M1021_g N_A_27_74#_c_484_n 5.80996e-19 $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_M1021_g N_A_27_74#_c_487_n 0.00746156f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_M1021_g N_A_27_74#_c_512_n 0.008978f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_c_210_n N_A_27_392#_c_675_n 7.39283e-19 $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_196 N_A_c_210_n N_A_27_392#_c_676_n 0.0122678f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_197 N_A_c_211_n N_A_27_392#_c_676_n 0.0126746f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_198 A N_A_27_392#_c_676_n 0.0246679f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_199 N_A_c_209_n N_A_27_392#_c_676_n 0.00372856f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_200 N_A_c_210_n N_A_116_392#_c_751_n 0.0124723f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_201 N_A_c_211_n N_A_116_392#_c_751_n 0.0147779f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_202 N_A_c_210_n N_A_116_392#_c_747_n 0.00447729f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_203 N_A_c_211_n N_A_116_392#_c_748_n 0.00283124f $X=1.405 $Y=1.885 $X2=0
+ $Y2=0
cc_204 N_A_c_210_n N_VPWR_c_771_n 0.00764661f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_205 N_A_c_211_n N_VPWR_c_771_n 0.00750914f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_206 N_A_c_210_n N_VPWR_c_776_n 0.00413917f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_207 N_A_c_211_n N_VPWR_c_777_n 0.00413917f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_208 N_A_c_210_n N_VPWR_c_770_n 0.0081781f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_209 N_A_c_211_n N_VPWR_c_770_n 0.00818241f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_210 N_A_M1021_g N_VGND_c_950_n 0.00478792f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_M1021_g N_VGND_c_957_n 0.00433162f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_M1021_g N_VGND_c_965_n 0.00437472f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_213 N_C_c_257_n N_A_563_48#_M1019_g 0.0048669f $X=3.935 $Y=1.295 $X2=0 $Y2=0
cc_214 N_C_c_258_n N_A_563_48#_M1019_g 0.00154557f $X=2.785 $Y=1.295 $X2=0 $Y2=0
cc_215 N_C_c_261_n N_A_563_48#_M1019_g 0.0178294f $X=2.41 $Y=1.385 $X2=0 $Y2=0
cc_216 N_C_c_262_n N_A_563_48#_M1019_g 0.0204994f $X=2.41 $Y=1.22 $X2=0 $Y2=0
cc_217 N_C_c_264_n N_A_563_48#_M1019_g 0.00457493f $X=2.64 $Y=1.295 $X2=0 $Y2=0
cc_218 N_C_c_266_n N_A_563_48#_c_356_n 0.0346776f $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_219 N_C_c_268_n N_A_563_48#_c_357_n 0.0363037f $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_220 N_C_c_257_n N_A_563_48#_c_351_n 0.00541921f $X=3.935 $Y=1.295 $X2=0 $Y2=0
cc_221 N_C_c_260_n N_A_563_48#_c_351_n 0.00179006f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_222 N_C_c_263_n N_A_563_48#_c_351_n 0.0169175f $X=4.03 $Y=1.345 $X2=0 $Y2=0
cc_223 N_C_c_263_n N_A_563_48#_c_352_n 9.5714e-19 $X=4.03 $Y=1.345 $X2=0 $Y2=0
cc_224 N_C_c_256_n N_A_563_48#_c_358_n 0.00683039f $X=3.805 $Y=1.795 $X2=0 $Y2=0
cc_225 N_C_c_268_n N_A_563_48#_c_358_n 0.00858865f $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_226 N_C_c_257_n N_A_563_48#_c_358_n 0.00801702f $X=3.935 $Y=1.295 $X2=0 $Y2=0
cc_227 N_C_c_259_n N_A_563_48#_c_358_n 0.00279021f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_228 N_C_c_260_n N_A_563_48#_c_358_n 0.0190105f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_229 N_C_c_263_n N_A_563_48#_c_358_n 0.00201502f $X=4.03 $Y=1.345 $X2=0 $Y2=0
cc_230 N_C_c_257_n N_A_563_48#_c_354_n 0.0122919f $X=3.935 $Y=1.295 $X2=0 $Y2=0
cc_231 N_C_c_260_n N_A_563_48#_c_354_n 0.00257448f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_232 N_C_c_263_n N_A_563_48#_c_354_n 0.00590433f $X=4.03 $Y=1.345 $X2=0 $Y2=0
cc_233 N_C_c_268_n N_A_563_48#_c_360_n 0.00551754f $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_234 N_C_c_255_n N_A_563_48#_c_355_n 0.0128898f $X=2.405 $Y=1.795 $X2=0 $Y2=0
cc_235 N_C_c_268_n N_A_563_48#_c_355_n 0.00360892f $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_236 N_C_c_257_n N_A_563_48#_c_355_n 0.00428911f $X=3.935 $Y=1.295 $X2=0 $Y2=0
cc_237 N_C_c_263_n N_A_563_48#_c_355_n 0.0201846f $X=4.03 $Y=1.345 $X2=0 $Y2=0
cc_238 N_C_c_263_n N_D_N_c_444_n 0.00113562f $X=4.03 $Y=1.345 $X2=-0.19
+ $Y2=-0.245
cc_239 N_C_c_256_n N_D_N_c_445_n 5.86466e-19 $X=3.805 $Y=1.795 $X2=0 $Y2=0
cc_240 N_C_c_260_n N_D_N_c_445_n 4.80178e-19 $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_241 N_C_c_263_n N_D_N_c_445_n 0.0132029f $X=4.03 $Y=1.345 $X2=0 $Y2=0
cc_242 N_C_c_256_n D_N 6.90614e-19 $X=3.805 $Y=1.795 $X2=0 $Y2=0
cc_243 N_C_c_259_n D_N 0.00725309f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_244 N_C_c_260_n D_N 0.0160858f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_245 N_C_c_263_n D_N 0.00207219f $X=4.03 $Y=1.345 $X2=0 $Y2=0
cc_246 N_C_c_257_n N_A_27_74#_c_488_n 0.0146246f $X=3.935 $Y=1.295 $X2=0 $Y2=0
cc_247 N_C_c_258_n N_A_27_74#_c_488_n 0.00874552f $X=2.785 $Y=1.295 $X2=0 $Y2=0
cc_248 N_C_c_261_n N_A_27_74#_c_488_n 9.3306e-19 $X=2.41 $Y=1.385 $X2=0 $Y2=0
cc_249 N_C_c_262_n N_A_27_74#_c_488_n 0.0158504f $X=2.41 $Y=1.22 $X2=0 $Y2=0
cc_250 N_C_c_264_n N_A_27_74#_c_488_n 0.0240592f $X=2.64 $Y=1.295 $X2=0 $Y2=0
cc_251 N_C_c_262_n N_A_27_74#_c_489_n 6.12903e-19 $X=2.41 $Y=1.22 $X2=0 $Y2=0
cc_252 N_C_c_255_n N_A_27_74#_c_490_n 7.49226e-19 $X=2.405 $Y=1.795 $X2=0 $Y2=0
cc_253 N_C_c_266_n N_A_27_74#_c_490_n 5.77326e-19 $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_254 N_C_c_257_n N_A_27_74#_c_490_n 0.0263933f $X=3.935 $Y=1.295 $X2=0 $Y2=0
cc_255 N_C_c_258_n N_A_27_74#_c_490_n 0.00272529f $X=2.785 $Y=1.295 $X2=0 $Y2=0
cc_256 N_C_c_261_n N_A_27_74#_c_490_n 3.38032e-19 $X=2.41 $Y=1.385 $X2=0 $Y2=0
cc_257 N_C_c_264_n N_A_27_74#_c_490_n 0.0442277f $X=2.64 $Y=1.295 $X2=0 $Y2=0
cc_258 N_C_c_257_n N_A_27_74#_c_491_n 0.0193845f $X=3.935 $Y=1.295 $X2=0 $Y2=0
cc_259 N_C_c_259_n N_A_27_74#_c_491_n 0.00343689f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_260 N_C_c_260_n N_A_27_74#_c_491_n 0.0212279f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_261 N_C_c_263_n N_A_27_74#_c_491_n 0.00768642f $X=4.03 $Y=1.345 $X2=0 $Y2=0
cc_262 N_C_c_262_n N_A_27_74#_c_494_n 0.00819477f $X=2.41 $Y=1.22 $X2=0 $Y2=0
cc_263 N_C_c_266_n N_A_27_74#_c_534_n 5.68706e-19 $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_264 N_C_c_268_n N_A_27_74#_c_534_n 5.77365e-19 $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_265 N_C_c_266_n N_A_27_392#_c_677_n 0.00376379f $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_266 N_C_c_261_n N_A_27_392#_c_677_n 3.26748e-19 $X=2.41 $Y=1.385 $X2=0 $Y2=0
cc_267 N_C_c_264_n N_A_27_392#_c_677_n 0.00903914f $X=2.64 $Y=1.295 $X2=0 $Y2=0
cc_268 N_C_c_266_n N_A_27_392#_c_702_n 0.00434089f $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_269 N_C_c_266_n N_A_27_392#_c_678_n 0.00617104f $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_270 N_C_c_266_n N_A_27_392#_c_704_n 0.0110243f $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_271 N_C_c_268_n N_A_27_392#_c_704_n 0.0134276f $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_272 N_C_c_264_n N_A_27_392#_c_704_n 0.0110956f $X=2.64 $Y=1.295 $X2=0 $Y2=0
cc_273 N_C_c_268_n N_A_27_392#_c_680_n 0.00667149f $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_274 N_C_c_266_n N_A_27_392#_c_708_n 2.24111e-19 $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_275 N_C_c_266_n N_VPWR_c_777_n 0.00445602f $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_276 N_C_c_268_n N_VPWR_c_777_n 0.00444483f $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_277 N_C_c_266_n N_VPWR_c_770_n 0.00445519f $X=2.405 $Y=1.885 $X2=0 $Y2=0
cc_278 N_C_c_268_n N_VPWR_c_770_n 0.00450333f $X=3.805 $Y=1.885 $X2=0 $Y2=0
cc_279 N_C_c_266_n N_A_496_392#_c_860_n 0.00155487f $X=2.405 $Y=1.885 $X2=0
+ $Y2=0
cc_280 N_C_c_268_n N_A_496_392#_c_860_n 0.00356698f $X=3.805 $Y=1.885 $X2=0
+ $Y2=0
cc_281 N_C_c_262_n N_VGND_c_951_n 0.00999028f $X=2.41 $Y=1.22 $X2=0 $Y2=0
cc_282 N_C_c_262_n N_VGND_c_957_n 0.00383152f $X=2.41 $Y=1.22 $X2=0 $Y2=0
cc_283 N_C_c_262_n N_VGND_c_965_n 0.00374269f $X=2.41 $Y=1.22 $X2=0 $Y2=0
cc_284 N_A_563_48#_c_353_n N_D_N_c_444_n 0.00701529f $X=4.4 $Y=0.505 $X2=-0.19
+ $Y2=-0.245
cc_285 N_A_563_48#_c_358_n N_D_N_c_445_n 0.00840209f $X=4.425 $Y=1.805 $X2=0
+ $Y2=0
cc_286 N_A_563_48#_c_360_n N_D_N_c_445_n 0.0106589f $X=4.59 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A_563_48#_c_358_n D_N 0.0264202f $X=4.425 $Y=1.805 $X2=0 $Y2=0
cc_288 N_A_563_48#_c_358_n N_A_27_74#_c_496_n 2.61985e-19 $X=4.425 $Y=1.805
+ $X2=0 $Y2=0
cc_289 N_A_563_48#_M1019_g N_A_27_74#_c_488_n 0.0141605f $X=2.89 $Y=0.74 $X2=0
+ $Y2=0
cc_290 N_A_563_48#_c_351_n N_A_27_74#_c_488_n 0.00796185f $X=3.4 $Y=1.47 $X2=0
+ $Y2=0
cc_291 N_A_563_48#_c_354_n N_A_27_74#_c_488_n 9.33451e-19 $X=3.635 $Y=1.805
+ $X2=0 $Y2=0
cc_292 N_A_563_48#_c_355_n N_A_27_74#_c_488_n 0.00630411f $X=3.355 $Y=1.677
+ $X2=0 $Y2=0
cc_293 N_A_563_48#_M1019_g N_A_27_74#_c_489_n 0.00901529f $X=2.89 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_563_48#_c_352_n N_A_27_74#_c_489_n 0.00406215f $X=3.605 $Y=0.505
+ $X2=0 $Y2=0
cc_295 N_A_563_48#_c_353_n N_A_27_74#_c_489_n 0.0270256f $X=4.4 $Y=0.505 $X2=0
+ $Y2=0
cc_296 N_A_563_48#_M1019_g N_A_27_74#_c_490_n 0.0070275f $X=2.89 $Y=0.74 $X2=0
+ $Y2=0
cc_297 N_A_563_48#_c_356_n N_A_27_74#_c_490_n 0.00367822f $X=2.905 $Y=1.885
+ $X2=0 $Y2=0
cc_298 N_A_563_48#_c_357_n N_A_27_74#_c_490_n 0.00241007f $X=3.355 $Y=1.885
+ $X2=0 $Y2=0
cc_299 N_A_563_48#_c_351_n N_A_27_74#_c_490_n 0.00583124f $X=3.4 $Y=1.47 $X2=0
+ $Y2=0
cc_300 N_A_563_48#_c_354_n N_A_27_74#_c_490_n 0.0284993f $X=3.635 $Y=1.805 $X2=0
+ $Y2=0
cc_301 N_A_563_48#_c_355_n N_A_27_74#_c_490_n 0.0168658f $X=3.355 $Y=1.677 $X2=0
+ $Y2=0
cc_302 N_A_563_48#_M1016_s N_A_27_74#_c_491_n 0.00665269f $X=3.88 $Y=0.36 $X2=0
+ $Y2=0
cc_303 N_A_563_48#_c_351_n N_A_27_74#_c_491_n 0.0138798f $X=3.4 $Y=1.47 $X2=0
+ $Y2=0
cc_304 N_A_563_48#_c_352_n N_A_27_74#_c_491_n 0.00586918f $X=3.605 $Y=0.505
+ $X2=0 $Y2=0
cc_305 N_A_563_48#_c_353_n N_A_27_74#_c_491_n 0.0829706f $X=4.4 $Y=0.505 $X2=0
+ $Y2=0
cc_306 N_A_563_48#_c_354_n N_A_27_74#_c_491_n 0.00605079f $X=3.635 $Y=1.805
+ $X2=0 $Y2=0
cc_307 N_A_563_48#_c_356_n N_A_27_74#_c_534_n 0.00511774f $X=2.905 $Y=1.885
+ $X2=0 $Y2=0
cc_308 N_A_563_48#_c_357_n N_A_27_74#_c_534_n 0.00354462f $X=3.355 $Y=1.885
+ $X2=0 $Y2=0
cc_309 N_A_563_48#_c_354_n N_A_27_74#_c_534_n 0.00222783f $X=3.635 $Y=1.805
+ $X2=0 $Y2=0
cc_310 N_A_563_48#_c_355_n N_A_27_74#_c_534_n 0.0061731f $X=3.355 $Y=1.677 $X2=0
+ $Y2=0
cc_311 N_A_563_48#_c_358_n N_A_27_74#_c_495_n 2.05886e-19 $X=4.425 $Y=1.805
+ $X2=0 $Y2=0
cc_312 N_A_563_48#_c_356_n N_A_27_392#_c_677_n 5.04162e-19 $X=2.905 $Y=1.885
+ $X2=0 $Y2=0
cc_313 N_A_563_48#_c_356_n N_A_27_392#_c_702_n 9.95667e-19 $X=2.905 $Y=1.885
+ $X2=0 $Y2=0
cc_314 N_A_563_48#_c_356_n N_A_27_392#_c_678_n 6.4283e-19 $X=2.905 $Y=1.885
+ $X2=0 $Y2=0
cc_315 N_A_563_48#_c_356_n N_A_27_392#_c_704_n 0.0129089f $X=2.905 $Y=1.885
+ $X2=0 $Y2=0
cc_316 N_A_563_48#_c_357_n N_A_27_392#_c_704_n 0.0123757f $X=3.355 $Y=1.885
+ $X2=0 $Y2=0
cc_317 N_A_563_48#_c_358_n N_A_27_392#_c_704_n 0.00817137f $X=4.425 $Y=1.805
+ $X2=0 $Y2=0
cc_318 N_A_563_48#_c_354_n N_A_27_392#_c_704_n 0.0103012f $X=3.635 $Y=1.805
+ $X2=0 $Y2=0
cc_319 N_A_563_48#_c_358_n N_A_27_392#_c_679_n 0.0205407f $X=4.425 $Y=1.805
+ $X2=0 $Y2=0
cc_320 N_A_563_48#_c_360_n N_A_27_392#_c_679_n 0.019777f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_321 N_A_563_48#_c_360_n N_A_27_392#_c_680_n 0.0217579f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_A_563_48#_c_360_n N_A_27_392#_c_681_n 0.0121617f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_563_48#_c_358_n N_VPWR_c_772_n 0.00491877f $X=4.425 $Y=1.805 $X2=0
+ $Y2=0
cc_324 N_A_563_48#_c_360_n N_VPWR_c_772_n 0.0638161f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A_563_48#_c_356_n N_VPWR_c_777_n 0.00291649f $X=2.905 $Y=1.885 $X2=0
+ $Y2=0
cc_326 N_A_563_48#_c_357_n N_VPWR_c_777_n 0.00291649f $X=3.355 $Y=1.885 $X2=0
+ $Y2=0
cc_327 N_A_563_48#_c_360_n N_VPWR_c_777_n 0.0097982f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_328 N_A_563_48#_c_356_n N_VPWR_c_770_n 0.0036003f $X=2.905 $Y=1.885 $X2=0
+ $Y2=0
cc_329 N_A_563_48#_c_357_n N_VPWR_c_770_n 0.00359599f $X=3.355 $Y=1.885 $X2=0
+ $Y2=0
cc_330 N_A_563_48#_c_360_n N_VPWR_c_770_n 0.0111907f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_331 N_A_563_48#_c_356_n N_A_496_392#_c_860_n 0.0111962f $X=2.905 $Y=1.885
+ $X2=0 $Y2=0
cc_332 N_A_563_48#_c_357_n N_A_496_392#_c_860_n 0.0112134f $X=3.355 $Y=1.885
+ $X2=0 $Y2=0
cc_333 N_A_563_48#_M1019_g N_VGND_c_951_n 0.00519744f $X=2.89 $Y=0.74 $X2=0
+ $Y2=0
cc_334 N_A_563_48#_c_353_n N_VGND_c_952_n 0.00839618f $X=4.4 $Y=0.505 $X2=0
+ $Y2=0
cc_335 N_A_563_48#_M1019_g N_VGND_c_958_n 0.00383287f $X=2.89 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A_563_48#_c_352_n N_VGND_c_958_n 0.0107668f $X=3.605 $Y=0.505 $X2=0
+ $Y2=0
cc_337 N_A_563_48#_c_353_n N_VGND_c_958_n 0.0485352f $X=4.4 $Y=0.505 $X2=0 $Y2=0
cc_338 N_A_563_48#_M1019_g N_VGND_c_965_n 0.00411093f $X=2.89 $Y=0.74 $X2=0
+ $Y2=0
cc_339 N_A_563_48#_c_352_n N_VGND_c_965_n 0.0141143f $X=3.605 $Y=0.505 $X2=0
+ $Y2=0
cc_340 N_A_563_48#_c_353_n N_VGND_c_965_n 0.0405648f $X=4.4 $Y=0.505 $X2=0 $Y2=0
cc_341 N_D_N_c_444_n N_A_27_74#_M1001_g 0.0195674f $X=4.695 $Y=1.22 $X2=0 $Y2=0
cc_342 N_D_N_c_445_n N_A_27_74#_M1001_g 0.0224913f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_343 D_N N_A_27_74#_M1001_g 3.77003e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_344 N_D_N_c_445_n N_A_27_74#_c_496_n 0.0152047f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_345 N_D_N_c_444_n N_A_27_74#_c_491_n 0.0143342f $X=4.695 $Y=1.22 $X2=0 $Y2=0
cc_346 N_D_N_c_445_n N_A_27_74#_c_491_n 0.00411665f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_347 D_N N_A_27_74#_c_491_n 0.024416f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_348 N_D_N_c_444_n N_A_27_74#_c_492_n 0.00358702f $X=4.695 $Y=1.22 $X2=0 $Y2=0
cc_349 N_D_N_c_445_n N_A_27_74#_c_492_n 7.01612e-19 $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_350 D_N N_A_27_74#_c_492_n 0.0107433f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_351 N_D_N_c_445_n N_A_27_74#_c_493_n 0.00489004f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_352 D_N N_A_27_74#_c_493_n 0.0195474f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_353 N_D_N_c_445_n N_A_27_74#_c_495_n 0.00461336f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_354 N_D_N_c_445_n N_A_27_392#_c_680_n 0.00323587f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_D_N_c_445_n N_VPWR_c_772_n 0.0121288f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_356 N_D_N_c_445_n N_VPWR_c_777_n 0.00481995f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_357 N_D_N_c_445_n N_VPWR_c_770_n 0.00508379f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_358 N_D_N_c_444_n N_VGND_c_952_n 0.00241507f $X=4.695 $Y=1.22 $X2=0 $Y2=0
cc_359 N_D_N_c_444_n N_VGND_c_958_n 0.00507111f $X=4.695 $Y=1.22 $X2=0 $Y2=0
cc_360 N_D_N_c_444_n N_VGND_c_965_n 0.00514438f $X=4.695 $Y=1.22 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_490_n N_A_27_392#_c_677_n 0.00202659f $X=2.98 $Y=2.02 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_534_n N_A_27_392#_c_677_n 0.00305196f $X=3.13 $Y=2.105 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_534_n N_A_27_392#_c_702_n 0.0019933f $X=3.13 $Y=2.105 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_M1008_d N_A_27_392#_c_704_n 0.00374176f $X=2.98 $Y=1.96 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_c_534_n N_A_27_392#_c_704_n 0.0201862f $X=3.13 $Y=2.105 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_534_n N_A_27_392#_c_679_n 0.0034257f $X=3.13 $Y=2.105 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_496_n N_VPWR_c_772_n 0.00769626f $X=5.35 $Y=1.765 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_493_n N_VPWR_c_772_n 0.0158832f $X=5.155 $Y=1.485 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_581_p N_VPWR_c_772_n 0.0045163f $X=5.99 $Y=1.485 $X2=0 $Y2=0
cc_370 N_A_27_74#_c_495_n N_VPWR_c_772_n 0.00154915f $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_496_n N_VPWR_c_773_n 5.28947e-19 $X=5.35 $Y=1.765 $X2=0
+ $Y2=0
cc_372 N_A_27_74#_c_497_n N_VPWR_c_773_n 0.0106488f $X=5.8 $Y=1.765 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_498_n N_VPWR_c_773_n 0.0105176f $X=6.25 $Y=1.765 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_499_n N_VPWR_c_773_n 4.98648e-19 $X=6.7 $Y=1.765 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_498_n N_VPWR_c_775_n 4.98648e-19 $X=6.25 $Y=1.765 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_499_n N_VPWR_c_775_n 0.0116621f $X=6.7 $Y=1.765 $X2=0 $Y2=0
cc_377 N_A_27_74#_c_496_n N_VPWR_c_778_n 0.00445602f $X=5.35 $Y=1.765 $X2=0
+ $Y2=0
cc_378 N_A_27_74#_c_497_n N_VPWR_c_778_n 0.00413917f $X=5.8 $Y=1.765 $X2=0 $Y2=0
cc_379 N_A_27_74#_c_498_n N_VPWR_c_779_n 0.00413917f $X=6.25 $Y=1.765 $X2=0
+ $Y2=0
cc_380 N_A_27_74#_c_499_n N_VPWR_c_779_n 0.00413917f $X=6.7 $Y=1.765 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_496_n N_VPWR_c_770_n 0.00862391f $X=5.35 $Y=1.765 $X2=0
+ $Y2=0
cc_382 N_A_27_74#_c_497_n N_VPWR_c_770_n 0.00817726f $X=5.8 $Y=1.765 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_498_n N_VPWR_c_770_n 0.00817726f $X=6.25 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_c_499_n N_VPWR_c_770_n 0.00817726f $X=6.7 $Y=1.765 $X2=0 $Y2=0
cc_385 N_A_27_74#_M1008_d N_A_496_392#_c_860_n 0.00201274f $X=2.98 $Y=1.96 $X2=0
+ $Y2=0
cc_386 N_A_27_74#_M1001_g N_X_c_873_n 5.50956e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_387 N_A_27_74#_M1013_g N_X_c_873_n 0.00377577f $X=5.775 $Y=0.74 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_496_n N_X_c_880_n 0.00387231f $X=5.35 $Y=1.765 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_581_p N_X_c_880_n 0.0235455f $X=5.99 $Y=1.485 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_495_n N_X_c_880_n 0.00656597f $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_391 N_A_27_74#_c_496_n N_X_c_881_n 0.00939243f $X=5.35 $Y=1.765 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_497_n N_X_c_881_n 3.88029e-19 $X=5.8 $Y=1.765 $X2=0 $Y2=0
cc_393 N_A_27_74#_M1013_g N_X_c_874_n 0.015091f $X=5.775 $Y=0.74 $X2=0 $Y2=0
cc_394 N_A_27_74#_M1014_g N_X_c_874_n 0.0133712f $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_395 N_A_27_74#_c_581_p N_X_c_874_n 0.036982f $X=5.99 $Y=1.485 $X2=0 $Y2=0
cc_396 N_A_27_74#_c_495_n N_X_c_874_n 0.00381149f $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_397 N_A_27_74#_M1001_g N_X_c_875_n 4.02336e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_398 N_A_27_74#_c_492_n N_X_c_875_n 0.00655124f $X=5.07 $Y=1.32 $X2=0 $Y2=0
cc_399 N_A_27_74#_c_581_p N_X_c_875_n 0.0278321f $X=5.99 $Y=1.485 $X2=0 $Y2=0
cc_400 N_A_27_74#_c_495_n N_X_c_875_n 0.00542073f $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_401 N_A_27_74#_c_497_n N_X_c_882_n 0.0177404f $X=5.8 $Y=1.765 $X2=0 $Y2=0
cc_402 N_A_27_74#_c_498_n N_X_c_882_n 0.0198915f $X=6.25 $Y=1.765 $X2=0 $Y2=0
cc_403 N_A_27_74#_c_581_p N_X_c_882_n 0.0361437f $X=5.99 $Y=1.485 $X2=0 $Y2=0
cc_404 N_A_27_74#_c_495_n N_X_c_882_n 0.00967485f $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_405 N_A_27_74#_M1013_g N_X_c_876_n 6.75677e-19 $X=5.775 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A_27_74#_M1014_g N_X_c_876_n 0.00903544f $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_407 N_A_27_74#_M1017_g N_X_c_876_n 3.97481e-19 $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_408 N_A_27_74#_c_498_n N_X_c_883_n 3.85296e-19 $X=6.25 $Y=1.765 $X2=0 $Y2=0
cc_409 N_A_27_74#_c_499_n N_X_c_883_n 3.85296e-19 $X=6.7 $Y=1.765 $X2=0 $Y2=0
cc_410 N_A_27_74#_c_498_n N_X_c_884_n 0.0014694f $X=6.25 $Y=1.765 $X2=0 $Y2=0
cc_411 N_A_27_74#_c_499_n N_X_c_884_n 0.00283006f $X=6.7 $Y=1.765 $X2=0 $Y2=0
cc_412 N_A_27_74#_c_581_p N_X_c_884_n 0.01197f $X=5.99 $Y=1.485 $X2=0 $Y2=0
cc_413 N_A_27_74#_c_495_n N_X_c_884_n 0.030378f $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_414 N_A_27_74#_M1014_g N_X_c_877_n 7.4184e-19 $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_415 N_A_27_74#_M1017_g N_X_c_877_n 7.94511e-19 $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_416 N_A_27_74#_M1013_g N_X_c_878_n 7.96351e-19 $X=5.775 $Y=0.74 $X2=0 $Y2=0
cc_417 N_A_27_74#_M1014_g N_X_c_878_n 0.0041295f $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_418 N_A_27_74#_M1017_g N_X_c_878_n 0.00381078f $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_419 N_A_27_74#_M1014_g N_X_c_879_n 5.95443e-19 $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_420 N_A_27_74#_M1017_g N_X_c_879_n 0.00229816f $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_421 N_A_27_74#_c_581_p N_X_c_879_n 0.0118939f $X=5.99 $Y=1.485 $X2=0 $Y2=0
cc_422 N_A_27_74#_c_495_n N_X_c_879_n 0.0159431f $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_423 N_A_27_74#_c_499_n X 0.00259717f $X=6.7 $Y=1.765 $X2=0 $Y2=0
cc_424 N_A_27_74#_c_499_n X 0.0211705f $X=6.7 $Y=1.765 $X2=0 $Y2=0
cc_425 N_A_27_74#_c_495_n X 7.03953e-19 $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_426 N_A_27_74#_c_512_n N_VGND_M1020_d 0.00692878f $X=1.115 $Y=0.645 $X2=-0.19
+ $Y2=-0.245
cc_427 N_A_27_74#_c_488_n N_VGND_M1018_d 0.00735178f $X=2.895 $Y=0.855 $X2=0
+ $Y2=0
cc_428 N_A_27_74#_c_491_n N_VGND_M1016_d 0.00685527f $X=4.985 $Y=0.925 $X2=0
+ $Y2=0
cc_429 N_A_27_74#_c_492_n N_VGND_M1016_d 0.00118596f $X=5.07 $Y=1.32 $X2=0 $Y2=0
cc_430 N_A_27_74#_c_484_n N_VGND_c_950_n 0.0101711f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_431 N_A_27_74#_c_487_n N_VGND_c_950_n 0.0112409f $X=1.41 $Y=0.645 $X2=0 $Y2=0
cc_432 N_A_27_74#_c_512_n N_VGND_c_950_n 0.0242009f $X=1.115 $Y=0.645 $X2=0
+ $Y2=0
cc_433 N_A_27_74#_c_488_n N_VGND_c_951_n 0.0227127f $X=2.895 $Y=0.855 $X2=0
+ $Y2=0
cc_434 N_A_27_74#_c_489_n N_VGND_c_951_n 0.0197319f $X=3.105 $Y=0.515 $X2=0
+ $Y2=0
cc_435 N_A_27_74#_c_494_n N_VGND_c_951_n 0.0103321f $X=2.2 $Y=0.645 $X2=0 $Y2=0
cc_436 N_A_27_74#_M1001_g N_VGND_c_952_n 0.00776616f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_437 N_A_27_74#_M1013_g N_VGND_c_952_n 3.99174e-19 $X=5.775 $Y=0.74 $X2=0
+ $Y2=0
cc_438 N_A_27_74#_c_491_n N_VGND_c_952_n 0.0223024f $X=4.985 $Y=0.925 $X2=0
+ $Y2=0
cc_439 N_A_27_74#_M1001_g N_VGND_c_953_n 4.39575e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_440 N_A_27_74#_M1013_g N_VGND_c_953_n 0.00995806f $X=5.775 $Y=0.74 $X2=0
+ $Y2=0
cc_441 N_A_27_74#_M1014_g N_VGND_c_953_n 0.00408259f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_442 N_A_27_74#_M1014_g N_VGND_c_955_n 6.13213e-19 $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_27_74#_M1017_g N_VGND_c_955_n 0.0160133f $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_444 N_A_27_74#_c_495_n N_VGND_c_955_n 3.66564e-19 $X=6.7 $Y=1.542 $X2=0 $Y2=0
cc_445 N_A_27_74#_c_484_n N_VGND_c_956_n 0.014415f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_446 N_A_27_74#_c_487_n N_VGND_c_957_n 0.0475979f $X=1.41 $Y=0.645 $X2=0 $Y2=0
cc_447 N_A_27_74#_c_489_n N_VGND_c_958_n 0.0164374f $X=3.105 $Y=0.515 $X2=0
+ $Y2=0
cc_448 N_A_27_74#_M1001_g N_VGND_c_959_n 0.00429299f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_449 N_A_27_74#_M1013_g N_VGND_c_959_n 0.00383152f $X=5.775 $Y=0.74 $X2=0
+ $Y2=0
cc_450 N_A_27_74#_M1014_g N_VGND_c_960_n 0.00434272f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_451 N_A_27_74#_M1017_g N_VGND_c_960_n 0.00383152f $X=6.705 $Y=0.74 $X2=0
+ $Y2=0
cc_452 N_A_27_74#_M1001_g N_VGND_c_965_n 0.0084864f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_453 N_A_27_74#_M1013_g N_VGND_c_965_n 0.00758657f $X=5.775 $Y=0.74 $X2=0
+ $Y2=0
cc_454 N_A_27_74#_M1014_g N_VGND_c_965_n 0.00820718f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_455 N_A_27_74#_M1017_g N_VGND_c_965_n 0.0075754f $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_456 N_A_27_74#_c_484_n N_VGND_c_965_n 0.0119404f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_457 N_A_27_74#_c_487_n N_VGND_c_965_n 0.0397185f $X=1.41 $Y=0.645 $X2=0 $Y2=0
cc_458 N_A_27_74#_c_488_n N_VGND_c_965_n 0.0123071f $X=2.895 $Y=0.855 $X2=0
+ $Y2=0
cc_459 N_A_27_74#_c_489_n N_VGND_c_965_n 0.0134433f $X=3.105 $Y=0.515 $X2=0
+ $Y2=0
cc_460 N_A_27_74#_c_491_n N_VGND_c_965_n 0.0166962f $X=4.985 $Y=0.925 $X2=0
+ $Y2=0
cc_461 N_A_27_74#_c_512_n N_VGND_c_965_n 0.0118956f $X=1.115 $Y=0.645 $X2=0
+ $Y2=0
cc_462 N_A_27_392#_c_676_n N_A_116_392#_M1006_d 0.00219763f $X=2.015 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_463 N_A_27_392#_c_676_n N_A_116_392#_M1010_s 0.00250873f $X=2.015 $Y=2.035
+ $X2=0 $Y2=0
cc_464 N_A_27_392#_c_676_n N_A_116_392#_c_751_n 0.0343548f $X=2.015 $Y=2.035
+ $X2=0 $Y2=0
cc_465 N_A_27_392#_c_675_n N_A_116_392#_c_747_n 0.046248f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_466 N_A_27_392#_c_676_n N_A_116_392#_c_747_n 0.0138473f $X=2.015 $Y=2.035
+ $X2=0 $Y2=0
cc_467 N_A_27_392#_c_676_n N_A_116_392#_c_748_n 0.0203253f $X=2.015 $Y=2.035
+ $X2=0 $Y2=0
cc_468 N_A_27_392#_c_678_n N_A_116_392#_c_748_n 0.0176756f $X=2.18 $Y=2.815
+ $X2=0 $Y2=0
cc_469 N_A_27_392#_c_676_n N_VPWR_M1007_d 0.00198204f $X=2.015 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_470 N_A_27_392#_c_675_n N_VPWR_c_776_n 0.0145938f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_471 N_A_27_392#_c_678_n N_VPWR_c_777_n 0.0145938f $X=2.18 $Y=2.815 $X2=0
+ $Y2=0
cc_472 N_A_27_392#_c_680_n N_VPWR_c_777_n 0.011066f $X=4.03 $Y=2.815 $X2=0 $Y2=0
cc_473 N_A_27_392#_c_675_n N_VPWR_c_770_n 0.0120466f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_474 N_A_27_392#_c_678_n N_VPWR_c_770_n 0.0120466f $X=2.18 $Y=2.815 $X2=0
+ $Y2=0
cc_475 N_A_27_392#_c_704_n N_VPWR_c_770_n 0.0130084f $X=3.945 $Y=2.445 $X2=0
+ $Y2=0
cc_476 N_A_27_392#_c_680_n N_VPWR_c_770_n 0.00915947f $X=4.03 $Y=2.815 $X2=0
+ $Y2=0
cc_477 N_A_27_392#_c_704_n N_A_496_392#_M1009_d 0.00797962f $X=3.945 $Y=2.445
+ $X2=-0.19 $Y2=1.66
cc_478 N_A_27_392#_c_704_n N_A_496_392#_M1012_s 0.00515422f $X=3.945 $Y=2.445
+ $X2=0 $Y2=0
cc_479 N_A_27_392#_c_678_n N_A_496_392#_c_860_n 0.0113199f $X=2.18 $Y=2.815
+ $X2=0 $Y2=0
cc_480 N_A_27_392#_c_704_n N_A_496_392#_c_860_n 0.0660711f $X=3.945 $Y=2.445
+ $X2=0 $Y2=0
cc_481 N_A_27_392#_c_680_n N_A_496_392#_c_860_n 0.0198191f $X=4.03 $Y=2.815
+ $X2=0 $Y2=0
cc_482 N_A_116_392#_c_751_n N_VPWR_M1007_d 0.00374424f $X=1.515 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_483 N_A_116_392#_c_751_n N_VPWR_c_771_n 0.0171814f $X=1.515 $Y=2.375 $X2=0
+ $Y2=0
cc_484 N_A_116_392#_c_747_n N_VPWR_c_771_n 0.0228252f $X=0.73 $Y=2.455 $X2=0
+ $Y2=0
cc_485 N_A_116_392#_c_748_n N_VPWR_c_771_n 0.0139233f $X=1.68 $Y=2.455 $X2=0
+ $Y2=0
cc_486 N_A_116_392#_c_747_n N_VPWR_c_776_n 0.00750433f $X=0.73 $Y=2.455 $X2=0
+ $Y2=0
cc_487 N_A_116_392#_c_748_n N_VPWR_c_777_n 0.0146094f $X=1.68 $Y=2.455 $X2=0
+ $Y2=0
cc_488 N_A_116_392#_c_747_n N_VPWR_c_770_n 0.00620791f $X=0.73 $Y=2.455 $X2=0
+ $Y2=0
cc_489 N_A_116_392#_c_748_n N_VPWR_c_770_n 0.0120527f $X=1.68 $Y=2.455 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_777_n N_A_496_392#_c_860_n 0.0504896f $X=4.96 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_770_n N_A_496_392#_c_860_n 0.0426127f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_772_n N_X_c_880_n 0.0235225f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_493 N_VPWR_c_772_n N_X_c_881_n 0.0549702f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_494 N_VPWR_c_773_n N_X_c_881_n 0.0255358f $X=6.025 $Y=2.405 $X2=0 $Y2=0
cc_495 N_VPWR_c_778_n N_X_c_881_n 0.0123628f $X=5.86 $Y=3.33 $X2=0 $Y2=0
cc_496 N_VPWR_c_770_n N_X_c_881_n 0.0101999f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_497 N_VPWR_M1002_s N_X_c_882_n 0.00201799f $X=5.875 $Y=1.84 $X2=0 $Y2=0
cc_498 N_VPWR_c_773_n N_X_c_882_n 0.0179913f $X=6.025 $Y=2.405 $X2=0 $Y2=0
cc_499 N_VPWR_c_773_n N_X_c_883_n 0.0255132f $X=6.025 $Y=2.405 $X2=0 $Y2=0
cc_500 N_VPWR_c_775_n N_X_c_883_n 0.0255132f $X=6.925 $Y=2.405 $X2=0 $Y2=0
cc_501 N_VPWR_c_779_n N_X_c_883_n 0.0101736f $X=6.76 $Y=3.33 $X2=0 $Y2=0
cc_502 N_VPWR_c_770_n N_X_c_883_n 0.0084208f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_503 N_VPWR_M1005_s X 0.00440927f $X=6.775 $Y=1.84 $X2=0 $Y2=0
cc_504 N_VPWR_c_775_n X 0.0218032f $X=6.925 $Y=2.405 $X2=0 $Y2=0
cc_505 N_X_c_874_n N_VGND_M1013_d 0.00250873f $X=6.325 $Y=1.065 $X2=0 $Y2=0
cc_506 N_X_c_873_n N_VGND_c_952_n 0.0127976f $X=5.49 $Y=0.515 $X2=0 $Y2=0
cc_507 N_X_c_873_n N_VGND_c_953_n 0.0180508f $X=5.49 $Y=0.515 $X2=0 $Y2=0
cc_508 N_X_c_874_n N_VGND_c_953_n 0.0210288f $X=6.325 $Y=1.065 $X2=0 $Y2=0
cc_509 N_X_c_876_n N_VGND_c_953_n 0.0173318f $X=6.49 $Y=0.515 $X2=0 $Y2=0
cc_510 N_X_c_876_n N_VGND_c_955_n 0.023308f $X=6.49 $Y=0.515 $X2=0 $Y2=0
cc_511 N_X_c_877_n N_VGND_c_955_n 0.00625076f $X=6.45 $Y=1.065 $X2=0 $Y2=0
cc_512 N_X_c_873_n N_VGND_c_959_n 0.0146357f $X=5.49 $Y=0.515 $X2=0 $Y2=0
cc_513 N_X_c_876_n N_VGND_c_960_n 0.0109942f $X=6.49 $Y=0.515 $X2=0 $Y2=0
cc_514 N_X_c_873_n N_VGND_c_965_n 0.0121141f $X=5.49 $Y=0.515 $X2=0 $Y2=0
cc_515 N_X_c_876_n N_VGND_c_965_n 0.00904371f $X=6.49 $Y=0.515 $X2=0 $Y2=0
