* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
M1000 a_664_392# a_231_74# a_586_392# VPB pshort w=1e+06u l=150000u
+  ad=3.278e+11p pd=2.76e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR a_863_98# a_770_508# VPB pshort w=420000u l=150000u
+  ad=2.07525e+12p pd=1.551e+07u as=2.121e+11p ps=1.85e+06u
M1002 VPWR a_863_98# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1003 a_231_74# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.4685e+12p ps=1.184e+07u
M1004 a_815_124# a_231_74# a_664_392# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.028e+11p ps=2.46e+06u
M1005 VPWR a_231_74# a_373_82# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1006 VGND D a_27_413# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1007 a_586_392# a_27_413# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_863_98# a_664_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1009 Q_N a_1347_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 a_770_508# a_373_82# a_664_392# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_863_98# a_664_392# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1012 a_664_392# a_373_82# a_589_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1013 a_589_80# a_27_413# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q_N a_1347_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.248e+11p pd=2.82e+06u as=0p ps=0u
M1015 VGND a_863_98# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1016 a_1347_424# a_863_98# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1017 VGND a_231_74# a_373_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1018 VPWR D a_27_413# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.436e+11p ps=2.26e+06u
M1019 VGND a_863_98# a_815_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_231_74# GATE VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1021 a_1347_424# a_863_98# VPWR VPB pshort w=840000u l=150000u
+  ad=2.436e+11p pd=2.26e+06u as=0p ps=0u
.ends
