* File: sky130_fd_sc_hs__and3_4.spice
* Created: Thu Aug 27 20:32:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__and3_4.pex.spice"
.subckt sky130_fd_sc_hs__and3_4  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_83_260#_M1007_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_83_260#_M1014_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1014_d N_A_83_260#_M1017_g N_X_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_83_260#_M1018_g N_X_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.133522 AS=0.1036 PD=1.16899 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1003 N_A_489_74#_M1003_d N_C_M1003_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.115478 PD=0.92 PS=1.01101 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1013 N_A_489_74#_M1003_d N_C_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_A_686_74#_M1000_d N_B_M1000_g N_A_489_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1024 PD=1.85 PS=0.96 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1001 N_A_686_74#_M1001_d N_B_M1001_g N_A_489_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=7.488 M=1 R=4.26667
+ SA=75000.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1005 N_A_83_260#_M1005_d N_A_M1005_g N_A_686_74#_M1001_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1184 AS=0.0896 PD=1.01 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1019 N_A_83_260#_M1005_d N_A_M1019_g N_A_686_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1184 AS=0.2144 PD=1.01 PS=1.95 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75001.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1006 N_X_M1006_d N_A_83_260#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75004.1 A=0.168 P=2.54 MULT=1
MM1008 N_X_M1006_d N_A_83_260#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75003.7 A=0.168 P=2.54 MULT=1
MM1009 N_X_M1009_d N_A_83_260#_M1009_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1009_d N_A_83_260#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2344 PD=1.42 PS=1.73714 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.7 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1011 N_A_83_260#_M1011_d N_C_M1011_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.1758 PD=1.14 PS=1.30286 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75002.2 SB=75003 A=0.126 P=1.98 MULT=1
MM1012 N_A_83_260#_M1011_d N_C_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.273 PD=1.14 PS=1.49 NRD=2.3443 NRS=3.5066 M=1 R=5.6 SA=75002.7
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1012_s N_B_M1004_g N_A_83_260#_M1004_s VPB PSHORT L=0.15 W=0.84
+ AD=0.273 AS=0.1428 PD=1.49 PS=1.18 NRD=3.5066 NRS=2.3443 M=1 R=5.6 SA=75003.5
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_B_M1016_g N_A_83_260#_M1004_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1428 PD=1.2 PS=1.18 NRD=4.6886 NRS=11.7215 M=1 R=5.6 SA=75004
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1016_d N_A_M1002_g N_A_83_260#_M1002_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.126 PD=1.2 PS=1.14 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75004.5
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_83_260#_M1002_s VPB PSHORT L=0.15 W=0.84
+ AD=0.2898 AS=0.126 PD=2.37 PS=1.14 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75004.9
+ SB=75000.3 A=0.126 P=1.98 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
c_53 VNB 0 1.52826e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__and3_4.pxi.spice"
*
.ends
*
*
