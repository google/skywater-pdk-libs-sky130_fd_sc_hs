* File: sky130_fd_sc_hs__a22o_4.pex.spice
* Created: Thu Aug 27 20:27:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A22O_4%A_95_306# 1 2 3 4 13 15 16 18 20 21 25 27 29
+ 30 31 32 34 35 37 38 40 41 43 44 46 50 52 53 55 60 67 70 71 74 75 77 78
c192 53 0 1.7358e-19 $X=2.56 $Y=2.905
c193 52 0 3.05957e-20 $X=2.56 $Y=1.68
c194 41 0 1.44963e-19 $X=2.645 $Y=1.35
r195 81 82 41.913 $w=3.45e-07 $l=3e-07 $layer=POLY_cond $X=1.915 $Y=1.557
+ $X2=2.215 $Y2=1.557
r196 80 81 18.1623 $w=3.45e-07 $l=1.3e-07 $layer=POLY_cond $X=1.785 $Y=1.557
+ $X2=1.915 $Y2=1.557
r197 77 78 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=1.145
+ $X2=5.725 $Y2=1.145
r198 75 78 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=3.96 $Y=1.18
+ $X2=5.725 $Y2=1.18
r199 73 75 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=1.132
+ $X2=3.96 $Y2=1.132
r200 73 74 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=1.132
+ $X2=3.63 $Y2=1.132
r201 69 71 5.21567 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.35 $Y=2.867
+ $X2=3.515 $Y2=2.867
r202 69 70 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.35 $Y=2.867
+ $X2=3.185 $Y2=2.867
r203 67 84 12.5739 $w=3.45e-07 $l=9e-08 $layer=POLY_cond $X=2.555 $Y=1.557
+ $X2=2.645 $Y2=1.557
r204 67 82 47.5014 $w=3.45e-07 $l=3.4e-07 $layer=POLY_cond $X=2.555 $Y=1.557
+ $X2=2.215 $Y2=1.557
r205 60 71 26.4702 $w=3.18e-07 $l=7.35e-07 $layer=LI1_cond $X=4.25 $Y=2.82
+ $X2=3.515 $Y2=2.82
r206 57 74 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.855 $Y=1.18
+ $X2=3.63 $Y2=1.18
r207 55 70 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.645 $Y=2.99
+ $X2=3.185 $Y2=2.99
r208 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=2.905
+ $X2=2.645 $Y2=2.99
r209 52 53 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=2.56 $Y=1.68
+ $X2=2.56 $Y2=2.905
r210 50 52 9.02084 $w=2.88e-07 $l=2.11069e-07 $layer=LI1_cond $X=2.665 $Y=1.515
+ $X2=2.56 $Y2=1.68
r211 50 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.555
+ $Y=1.515 $X2=2.555 $Y2=1.515
r212 50 57 14.191 $w=2.88e-07 $l=4.19375e-07 $layer=LI1_cond $X=2.665 $Y=1.515
+ $X2=2.855 $Y2=1.18
r213 48 49 25.8634 $w=2.05e-07 $l=1.1e-07 $layer=POLY_cond $X=1.355 $Y=1.647
+ $X2=1.465 $Y2=1.647
r214 41 84 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.645 $Y=1.35
+ $X2=2.645 $Y2=1.557
r215 41 43 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.645 $Y=1.35
+ $X2=2.645 $Y2=0.87
r216 38 82 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.215 $Y=1.35
+ $X2=2.215 $Y2=1.557
r217 38 40 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.215 $Y=1.35
+ $X2=2.215 $Y2=0.87
r218 35 81 22.2839 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.915 $Y=1.765
+ $X2=1.915 $Y2=1.557
r219 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.915 $Y=1.765
+ $X2=1.915 $Y2=2.4
r220 32 80 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.785 $Y=1.35
+ $X2=1.785 $Y2=1.557
r221 32 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.785 $Y=1.35
+ $X2=1.785 $Y2=0.87
r222 31 49 24.721 $w=2.05e-07 $l=1.08995e-07 $layer=POLY_cond $X=1.555 $Y=1.605
+ $X2=1.465 $Y2=1.647
r223 30 80 26.1549 $w=3.45e-07 $l=9.60469e-08 $layer=POLY_cond $X=1.71 $Y=1.605
+ $X2=1.785 $Y2=1.557
r224 30 31 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.71 $Y=1.605
+ $X2=1.555 $Y2=1.605
r225 27 49 10.146 $w=1.5e-07 $l=1.18e-07 $layer=POLY_cond $X=1.465 $Y=1.765
+ $X2=1.465 $Y2=1.647
r226 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.465 $Y=1.765
+ $X2=1.465 $Y2=2.4
r227 23 48 10.146 $w=1.5e-07 $l=1.17e-07 $layer=POLY_cond $X=1.355 $Y=1.53
+ $X2=1.355 $Y2=1.647
r228 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.355 $Y=1.53
+ $X2=1.355 $Y2=0.87
r229 22 46 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.105 $Y=1.605
+ $X2=1.015 $Y2=1.605
r230 21 48 21.1942 $w=2.05e-07 $l=9.3675e-08 $layer=POLY_cond $X=1.28 $Y=1.605
+ $X2=1.355 $Y2=1.647
r231 21 22 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.28 $Y=1.605
+ $X2=1.105 $Y2=1.605
r232 18 46 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=1.015 $Y=1.765
+ $X2=1.015 $Y2=1.605
r233 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.015 $Y=1.765
+ $X2=1.015 $Y2=2.4
r234 17 44 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.655 $Y=1.605
+ $X2=0.565 $Y2=1.605
r235 16 46 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.925 $Y=1.605
+ $X2=1.015 $Y2=1.605
r236 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.925 $Y=1.605
+ $X2=0.655 $Y2=1.605
r237 13 44 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=0.565 $Y=1.765
+ $X2=0.565 $Y2=1.605
r238 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.565 $Y=1.765
+ $X2=0.565 $Y2=2.4
r239 4 60 600 $w=1.7e-07 $l=8.91852e-07 $layer=licon1_PDIFF $count=1 $X=4.1
+ $Y=1.96 $X2=4.25 $Y2=2.78
r240 3 69 600 $w=1.7e-07 $l=8.91852e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.96 $X2=3.35 $Y2=2.78
r241 2 77 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.75
+ $Y=0.615 $X2=5.89 $Y2=1.105
r242 1 73 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.655
+ $Y=0.6 $X2=3.795 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%B2 1 3 6 8 10 13 16 18 19 21 28 30 31 32 38
c96 30 0 1.7358e-19 $X=3.325 $Y=2.042
c97 13 0 1.65576e-20 $X=4.485 $Y=0.935
c98 8 0 1.69887e-19 $X=4.475 $Y=1.885
r99 32 38 3.07165 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=2.042
+ $X2=4.025 $Y2=2.042
r100 32 38 0.80403 $w=2.13e-07 $l=1.5e-08 $layer=LI1_cond $X=4.01 $Y=2.042
+ $X2=4.025 $Y2=2.042
r101 31 32 21.9768 $w=2.13e-07 $l=4.1e-07 $layer=LI1_cond $X=3.6 $Y=2.042
+ $X2=4.01 $Y2=2.042
r102 30 31 14.7406 $w=2.13e-07 $l=2.75e-07 $layer=LI1_cond $X=3.325 $Y=2.042
+ $X2=3.6 $Y2=2.042
r103 25 28 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.11 $Y=1.6
+ $X2=3.24 $Y2=1.6
r104 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.6 $X2=3.11 $Y2=1.6
r105 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.49
+ $Y=1.605 $X2=4.49 $Y2=1.605
r106 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.195 $Y=1.605
+ $X2=4.49 $Y2=1.605
r107 18 32 3.86667 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=4.11 $Y=1.935
+ $X2=4.11 $Y2=2.042
r108 17 19 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.11 $Y=1.77
+ $X2=4.195 $Y2=1.605
r109 17 18 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.11 $Y=1.77
+ $X2=4.11 $Y2=1.935
r110 16 30 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.24 $Y=1.935
+ $X2=3.325 $Y2=2.042
r111 15 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=1.765
+ $X2=3.24 $Y2=1.6
r112 15 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.24 $Y=1.765
+ $X2=3.24 $Y2=1.935
r113 11 22 38.6072 $w=2.91e-07 $l=1.67481e-07 $layer=POLY_cond $X=4.485 $Y=1.44
+ $X2=4.49 $Y2=1.605
r114 11 13 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.485 $Y=1.44
+ $X2=4.485 $Y2=0.935
r115 8 22 57.6553 $w=2.91e-07 $l=2.87402e-07 $layer=POLY_cond $X=4.475 $Y=1.885
+ $X2=4.49 $Y2=1.605
r116 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.475 $Y=1.885
+ $X2=4.475 $Y2=2.46
r117 4 26 38.6157 $w=2.9e-07 $l=1.83916e-07 $layer=POLY_cond $X=3.15 $Y=1.435
+ $X2=3.11 $Y2=1.6
r118 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.15 $Y=1.435
+ $X2=3.15 $Y2=0.92
r119 1 26 58.5605 $w=2.9e-07 $l=2.92404e-07 $layer=POLY_cond $X=3.125 $Y=1.885
+ $X2=3.11 $Y2=1.6
r120 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.125 $Y=1.885
+ $X2=3.125 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%B1 1 3 6 10 12 14 15 22
c54 15 0 2.17041e-19 $X=3.6 $Y=1.665
r55 22 23 1.81658 $w=3.98e-07 $l=1.5e-08 $layer=POLY_cond $X=4.01 $Y=1.66
+ $X2=4.025 $Y2=1.66
r56 20 22 42.3869 $w=3.98e-07 $l=3.5e-07 $layer=POLY_cond $X=3.66 $Y=1.66
+ $X2=4.01 $Y2=1.66
r57 18 20 9.68844 $w=3.98e-07 $l=8e-08 $layer=POLY_cond $X=3.58 $Y=1.66 $X2=3.66
+ $Y2=1.66
r58 17 18 0.605528 $w=3.98e-07 $l=5e-09 $layer=POLY_cond $X=3.575 $Y=1.66
+ $X2=3.58 $Y2=1.66
r59 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=1.6 $X2=3.66 $Y2=1.6
r60 12 23 25.7394 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.025 $Y=1.885
+ $X2=4.025 $Y2=1.66
r61 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.025 $Y=1.885
+ $X2=4.025 $Y2=2.46
r62 8 22 25.7394 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.01 $Y=1.435
+ $X2=4.01 $Y2=1.66
r63 8 10 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.01 $Y=1.435
+ $X2=4.01 $Y2=0.92
r64 4 18 25.7394 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=3.58 $Y=1.435
+ $X2=3.58 $Y2=1.66
r65 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.58 $Y=1.435
+ $X2=3.58 $Y2=0.92
r66 1 17 25.7394 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=3.575 $Y=1.885
+ $X2=3.575 $Y2=1.66
r67 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.575 $Y=1.885
+ $X2=3.575 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%A1 1 3 6 8 10 13 15 16 24
c53 13 0 1.56257e-19 $X=6.105 $Y=0.935
c54 6 0 1.25428e-19 $X=5.675 $Y=0.935
r55 24 25 4.34794 $w=3.88e-07 $l=3.5e-08 $layer=POLY_cond $X=6.07 $Y=1.667
+ $X2=6.105 $Y2=1.667
r56 22 24 46.5851 $w=3.88e-07 $l=3.75e-07 $layer=POLY_cond $X=5.695 $Y=1.667
+ $X2=6.07 $Y2=1.667
r57 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.695
+ $Y=1.615 $X2=5.695 $Y2=1.615
r58 20 22 2.48454 $w=3.88e-07 $l=2e-08 $layer=POLY_cond $X=5.675 $Y=1.667
+ $X2=5.695 $Y2=1.667
r59 19 20 6.83247 $w=3.88e-07 $l=5.5e-08 $layer=POLY_cond $X=5.62 $Y=1.667
+ $X2=5.675 $Y2=1.667
r60 16 23 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6 $Y=1.615
+ $X2=5.695 $Y2=1.615
r61 15 23 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=5.52 $Y=1.615
+ $X2=5.695 $Y2=1.615
r62 11 25 25.1189 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.105 $Y=1.45
+ $X2=6.105 $Y2=1.667
r63 11 13 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=6.105 $Y=1.45
+ $X2=6.105 $Y2=0.935
r64 8 24 25.1189 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.07 $Y=1.885
+ $X2=6.07 $Y2=1.667
r65 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.07 $Y=1.885
+ $X2=6.07 $Y2=2.46
r66 4 20 25.1189 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.675 $Y=1.45
+ $X2=5.675 $Y2=1.667
r67 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=5.675 $Y=1.45
+ $X2=5.675 $Y2=0.935
r68 1 19 25.1189 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.62 $Y=1.885
+ $X2=5.62 $Y2=1.667
r69 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.62 $Y=1.885
+ $X2=5.62 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%A2 2 3 5 9 10 12 13 14 16 20 23 26 28
c67 26 0 1.25428e-19 $X=5.04 $Y=0.555
c68 20 0 2.7975e-19 $X=6.535 $Y=0.935
c69 3 0 1.68376e-19 $X=4.955 $Y=1.885
r70 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=0.34
+ $X2=5.155 $Y2=0.505
r71 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=0.34 $X2=5.155 $Y2=0.34
r72 28 31 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.155 $Y=0.2
+ $X2=5.155 $Y2=0.34
r73 26 32 9.13937 $w=2.87e-07 $l=2.58998e-07 $layer=LI1_cond $X=5.04 $Y=0.555
+ $X2=5.137 $Y2=0.34
r74 20 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.535 $Y=0.935
+ $X2=6.535 $Y2=1.33
r75 17 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.535 $Y=0.275
+ $X2=6.535 $Y2=0.935
r76 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.52 $Y=1.885
+ $X2=6.52 $Y2=2.46
r77 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.52 $Y=1.795 $X2=6.52
+ $Y2=1.885
r78 12 25 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.52 $Y=1.42 $X2=6.52
+ $Y2=1.33
r79 12 13 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=6.52 $Y=1.42
+ $X2=6.52 $Y2=1.795
r80 11 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=0.2
+ $X2=5.155 $Y2=0.2
r81 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.46 $Y=0.2
+ $X2=6.535 $Y2=0.275
r82 10 11 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=6.46 $Y=0.2
+ $X2=5.32 $Y2=0.2
r83 9 33 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.245 $Y=0.935
+ $X2=5.245 $Y2=0.505
r84 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.245 $Y=1.33
+ $X2=5.245 $Y2=1.405
r85 7 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.245 $Y=1.33
+ $X2=5.245 $Y2=0.935
r86 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.955 $Y=1.885
+ $X2=4.955 $Y2=2.46
r87 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.955 $Y=1.795 $X2=4.955
+ $Y2=1.885
r88 1 23 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.955 $Y=1.405
+ $X2=5.245 $Y2=1.405
r89 1 2 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=4.955 $Y=1.48
+ $X2=4.955 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%VPWR 1 2 3 4 5 16 18 24 30 36 40 43 44 45 47
+ 52 57 67 68 74 77 80
r89 80 81 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r90 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r91 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r92 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r93 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r94 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r95 65 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r96 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r97 62 80 10.9443 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=5.51 $Y=3.33
+ $X2=5.272 $Y2=3.33
r98 62 64 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.51 $Y=3.33 $X2=6
+ $Y2=3.33
r99 61 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r100 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 58 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.18 $Y2=3.33
r102 58 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 57 80 10.9443 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.272 $Y2=3.33
r104 57 60 156.251 $w=1.68e-07 $l=2.395e-06 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 56 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 56 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 53 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 53 55 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 52 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.055 $Y=3.33
+ $X2=2.18 $Y2=3.33
r111 52 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.055 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 51 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r113 51 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r114 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 48 71 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.252 $Y2=3.33
r116 48 50 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 47 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 47 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 45 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 45 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r121 43 64 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.13 $Y=3.33 $X2=6
+ $Y2=3.33
r122 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.13 $Y=3.33
+ $X2=6.295 $Y2=3.33
r123 42 67 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.46 $Y=3.33 $X2=6.96
+ $Y2=3.33
r124 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.46 $Y=3.33
+ $X2=6.295 $Y2=3.33
r125 38 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=3.245
+ $X2=6.295 $Y2=3.33
r126 38 40 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.295 $Y=3.245
+ $X2=6.295 $Y2=2.375
r127 34 80 1.94084 $w=4.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.272 $Y=3.245
+ $X2=5.272 $Y2=3.33
r128 34 36 21.9071 $w=4.73e-07 $l=8.7e-07 $layer=LI1_cond $X=5.272 $Y=3.245
+ $X2=5.272 $Y2=2.375
r129 30 33 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=2.18 $Y=2.015
+ $X2=2.18 $Y2=2.815
r130 28 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=3.33
r131 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=2.815
r132 24 27 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.2 $Y2=2.815
r133 22 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=3.245
+ $X2=1.2 $Y2=3.33
r134 22 27 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=3.245 $X2=1.2
+ $Y2=2.815
r135 18 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.34 $Y=1.985
+ $X2=0.34 $Y2=2.815
r136 16 71 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.252 $Y2=3.33
r137 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.34 $Y2=2.815
r138 5 40 300 $w=1.7e-07 $l=4.84226e-07 $layer=licon1_PDIFF $count=2 $X=6.145
+ $Y=1.96 $X2=6.295 $Y2=2.375
r139 4 36 300 $w=1.7e-07 $l=5.21368e-07 $layer=licon1_PDIFF $count=2 $X=5.03
+ $Y=1.96 $X2=5.27 $Y2=2.375
r140 3 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.84 $X2=2.14 $Y2=2.815
r141 3 30 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.84 $X2=2.14 $Y2=2.015
r142 2 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.84 $X2=1.24 $Y2=2.815
r143 2 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.84 $X2=1.24 $Y2=1.985
r144 1 21 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.84 $X2=0.34 $Y2=2.815
r145 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.84 $X2=0.34 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%X 1 2 3 4 15 23 27 31 35 38 41 42 43 47
c67 35 0 1.44963e-19 $X=2.43 $Y=0.645
r68 43 47 2.47594 $w=3.9e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.79 $Y=1.395
+ $X2=0.705 $Y2=1.275
r69 43 47 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.67 $Y=1.275
+ $X2=0.705 $Y2=1.275
r70 42 43 18.3537 $w=2.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=1.275
+ $X2=0.67 $Y2=1.275
r71 40 41 10.4169 $w=6.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.69 $Y=1.33
+ $X2=1.855 $Y2=1.33
r72 39 40 2.9902 $w=6.38e-07 $l=1.6e-07 $layer=LI1_cond $X=1.53 $Y=1.33 $X2=1.69
+ $Y2=1.33
r73 38 39 2.86376 $w=6.38e-07 $l=1.25e-07 $layer=LI1_cond $X=1.405 $Y=1.33
+ $X2=1.53 $Y2=1.33
r74 33 35 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=2.39 $Y=1.01
+ $X2=2.39 $Y2=0.645
r75 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.265 $Y=1.095
+ $X2=2.39 $Y2=1.01
r76 31 41 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.265 $Y=1.095
+ $X2=1.855 $Y2=1.095
r77 27 29 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.69 $Y=1.985
+ $X2=1.69 $Y2=2.815
r78 25 40 4.6183 $w=3.3e-07 $l=3.2e-07 $layer=LI1_cond $X=1.69 $Y=1.65 $X2=1.69
+ $Y2=1.33
r79 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.69 $Y=1.65
+ $X2=1.69 $Y2=1.985
r80 21 39 6.29411 $w=2.5e-07 $l=3.2e-07 $layer=LI1_cond $X=1.53 $Y=1.01 $X2=1.53
+ $Y2=1.33
r81 21 23 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.53 $Y=1.01
+ $X2=1.53 $Y2=0.645
r82 20 43 2.47594 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=1.395
+ $X2=0.79 $Y2=1.395
r83 20 38 12.4298 $w=5.08e-07 $l=5.3e-07 $layer=LI1_cond $X=0.875 $Y=1.395
+ $X2=1.405 $Y2=1.395
r84 15 17 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=0.79 $Y=1.985
+ $X2=0.79 $Y2=2.815
r85 13 43 4.4465 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.79 $Y=1.65 $X2=0.79
+ $Y2=1.395
r86 13 15 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.79 $Y=1.65
+ $X2=0.79 $Y2=1.985
r87 4 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.84 $X2=1.69 $Y2=2.815
r88 4 27 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.84 $X2=1.69 $Y2=1.985
r89 3 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.84 $X2=0.79 $Y2=2.815
r90 3 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.84 $X2=0.79 $Y2=1.985
r91 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.5 $X2=2.43 $Y2=0.645
r92 1 39 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.5 $X2=1.57 $Y2=1.095
r93 1 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.5 $X2=1.57 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%A_555_392# 1 2 3 4 5 18 20 24 25 28 32 34 36
+ 38 40 47 49
c76 47 0 1.68376e-19 $X=4.7 $Y=2.46
r77 40 42 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=2.405
+ $X2=2.9 $Y2=2.57
r78 36 51 2.9222 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=6.785 $Y=2.12 $X2=6.785
+ $Y2=2.03
r79 36 38 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=6.785 $Y=2.12
+ $X2=6.785 $Y2=2.815
r80 35 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.93 $Y=2.035
+ $X2=5.805 $Y2=2.035
r81 34 51 4.22096 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=6.66 $Y=2.035
+ $X2=6.785 $Y2=2.03
r82 34 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.66 $Y=2.035
+ $X2=5.93 $Y2=2.035
r83 30 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.805 $Y=2.12
+ $X2=5.805 $Y2=2.035
r84 30 32 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.805 $Y=2.12
+ $X2=5.805 $Y2=2.815
r85 29 45 4.22096 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=4.865 $Y=2.035
+ $X2=4.74 $Y2=2.03
r86 28 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.68 $Y=2.035
+ $X2=5.805 $Y2=2.035
r87 28 29 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=5.68 $Y=2.035
+ $X2=4.865 $Y2=2.035
r88 25 47 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.74 $Y=2.32 $X2=4.74
+ $Y2=2.405
r89 24 45 2.9222 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=4.74 $Y=2.12 $X2=4.74
+ $Y2=2.03
r90 24 25 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=4.74 $Y=2.12 $X2=4.74
+ $Y2=2.32
r91 21 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=2.405
+ $X2=2.9 $Y2=2.405
r92 21 23 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.985 $Y=2.405
+ $X2=3.8 $Y2=2.405
r93 20 47 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.615 $Y=2.405
+ $X2=4.74 $Y2=2.405
r94 20 23 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=4.615 $Y=2.405
+ $X2=3.8 $Y2=2.405
r95 16 40 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=2.32 $X2=2.9
+ $Y2=2.405
r96 16 18 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.9 $Y=2.32 $X2=2.9
+ $Y2=2.105
r97 5 51 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.595
+ $Y=1.96 $X2=6.745 $Y2=2.105
r98 5 38 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.595
+ $Y=1.96 $X2=6.745 $Y2=2.815
r99 4 49 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=1.96 $X2=5.845 $Y2=2.115
r100 4 32 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=1.96 $X2=5.845 $Y2=2.815
r101 3 47 300 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_PDIFF $count=2 $X=4.55
+ $Y=1.96 $X2=4.7 $Y2=2.46
r102 3 45 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.55
+ $Y=1.96 $X2=4.7 $Y2=2.105
r103 2 23 600 $w=1.7e-07 $l=5.14563e-07 $layer=licon1_PDIFF $count=1 $X=3.65
+ $Y=1.96 $X2=3.8 $Y2=2.405
r104 1 42 600 $w=1.7e-07 $l=6.69589e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.96 $X2=2.9 $Y2=2.57
r105 1 18 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.96 $X2=2.9 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 45 46 47 48 60 73 75
r88 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r89 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r90 70 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r91 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r92 67 70 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r93 67 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r94 66 69 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r95 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r96 64 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=4.66
+ $Y2=0
r97 64 66 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=5.04
+ $Y2=0
r98 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r99 60 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.535 $Y=0 $X2=4.66
+ $Y2=0
r100 60 62 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=4.535 $Y=0
+ $X2=3.12 $Y2=0
r101 59 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r102 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r103 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r104 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r105 52 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r106 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r107 48 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r108 48 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r109 46 69 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.585 $Y=0
+ $X2=6.48 $Y2=0
r110 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=0 $X2=6.75
+ $Y2=0
r111 45 72 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.96
+ $Y2=0
r112 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.75
+ $Y2=0
r113 43 58 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.64
+ $Y2=0
r114 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.86
+ $Y2=0
r115 42 62 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.025 $Y=0 $X2=3.12
+ $Y2=0
r116 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=2.86
+ $Y2=0
r117 40 55 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=0
+ $X2=1.68 $Y2=0
r118 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.96
+ $Y2=0
r119 39 58 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.085 $Y=0
+ $X2=2.64 $Y2=0
r120 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=1.96
+ $Y2=0
r121 37 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r122 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.1
+ $Y2=0
r123 36 55 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.225 $Y=0
+ $X2=1.68 $Y2=0
r124 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.1
+ $Y2=0
r125 32 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.75 $Y=0.085
+ $X2=6.75 $Y2=0
r126 32 34 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.75 $Y=0.085
+ $X2=6.75 $Y2=0.76
r127 28 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0
r128 28 30 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0.76
r129 24 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0
r130 24 26 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0.75
r131 20 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r132 20 22 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.66
r133 16 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r134 16 18 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.805
r135 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.61
+ $Y=0.615 $X2=6.75 $Y2=0.76
r136 4 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.56
+ $Y=0.615 $X2=4.7 $Y2=0.76
r137 3 26 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.72
+ $Y=0.5 $X2=2.86 $Y2=0.75
r138 2 22 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.5 $X2=2 $Y2=0.66
r139 1 18 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.5 $X2=1.14 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%A_645_120# 1 2 12 13
r17 12 13 4.40113 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=4.245 $Y=0.752
+ $X2=4.14 $Y2=0.752
r18 9 13 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=3.365 $Y=0.705
+ $X2=4.14 $Y2=0.705
r19 2 12 182 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_NDIFF $count=1 $X=4.085
+ $Y=0.6 $X2=4.245 $Y2=0.75
r20 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.6 $X2=3.365 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_4%A_1064_123# 1 2 7 11 13
c23 13 0 2.96052e-19 $X=6.32 $Y=1.11
c24 11 0 1.39955e-19 $X=6.32 $Y=0.845
r25 11 16 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.32 $Y=0.845
+ $X2=6.32 $Y2=0.72
r26 11 13 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.32 $Y=0.845
+ $X2=6.32 $Y2=1.11
r27 7 16 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=6.235 $Y=0.76
+ $X2=6.32 $Y2=0.72
r28 7 9 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=6.235 $Y=0.76
+ $X2=5.46 $Y2=0.76
r29 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.18
+ $Y=0.615 $X2=6.32 $Y2=0.76
r30 2 13 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.18
+ $Y=0.615 $X2=6.32 $Y2=1.11
r31 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.615 $X2=5.46 $Y2=0.76
.ends

