* File: sky130_fd_sc_hs__dlxbn_2.pex.spice
* Created: Thu Aug 27 20:42:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DLXBN_2%D 3 6 7 9 10 13
c37 13 0 1.67694e-19 $X=0.605 $Y=1.615
c38 7 0 2.5702e-19 $X=0.59 $Y=2.045
r39 13 16 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.615
+ $X2=0.595 $Y2=1.78
r40 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.615
+ $X2=0.595 $Y2=1.45
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.615 $X2=0.605 $Y2=1.615
r42 10 14 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.605 $Y2=1.615
r43 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.59 $Y=2.045 $X2=0.59
+ $Y2=2.54
r44 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.59 $Y=1.955 $X2=0.59
+ $Y2=2.045
r45 6 16 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=0.59 $Y=1.955
+ $X2=0.59 $Y2=1.78
r46 3 15 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=0.955
+ $X2=0.495 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%GATE_N 3 5 7 8 12
c35 12 0 9.5906e-20 $X=1.15 $Y=1.795
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.795 $X2=1.15 $Y2=1.795
r37 8 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.15 $Y=2.035 $X2=1.15
+ $Y2=1.795
r38 5 11 52.2586 $w=2.99e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.09 $Y=2.045
+ $X2=1.15 $Y2=1.795
r39 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.09 $Y=2.045 $X2=1.09
+ $Y2=2.54
r40 1 11 38.5562 $w=2.99e-07 $l=1.94808e-07 $layer=POLY_cond $X=1.085 $Y=1.63
+ $X2=1.15 $Y2=1.795
r41 1 3 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.085 $Y=1.63 $X2=1.085
+ $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%A_232_98# 1 2 7 11 17 18 20 21 22 24 25 27
+ 28 29 30 33 35 38 39 42 47 55 60 62 67
c146 67 0 3.16539e-20 $X=3.995 $Y=1.652
c147 60 0 1.87089e-19 $X=4.19 $Y=1.585
c148 47 0 7.17879e-20 $X=1.72 $Y=1.425
c149 35 0 1.1467e-19 $X=1.317 $Y=2.56
c150 18 0 1.8903e-19 $X=3.16 $Y=1.11
r151 66 67 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=3.73 $Y=1.652
+ $X2=3.995 $Y2=1.652
r152 58 67 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=4.06 $Y=1.652
+ $X2=3.995 $Y2=1.652
r153 57 60 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.06 $Y=1.585
+ $X2=4.19 $Y2=1.585
r154 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=1.585 $X2=4.06 $Y2=1.585
r155 54 55 5.07737 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.44
+ $X2=1.655 $Y2=2.44
r156 48 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.72 $Y=1.425
+ $X2=1.72 $Y2=1.335
r157 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.425 $X2=1.72 $Y2=1.425
r158 45 47 6.52326 $w=2.63e-07 $l=1.5e-07 $layer=LI1_cond $X=1.57 $Y=1.392
+ $X2=1.72 $Y2=1.392
r159 41 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.19 $Y=1.75
+ $X2=4.19 $Y2=1.585
r160 41 42 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.19 $Y=1.75
+ $X2=4.19 $Y2=2.39
r161 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=2.475
+ $X2=4.19 $Y2=2.39
r162 39 55 159.84 $w=1.68e-07 $l=2.45e-06 $layer=LI1_cond $X=4.105 $Y=2.475
+ $X2=1.655 $Y2=2.475
r163 38 54 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.57 $Y=2.32
+ $X2=1.57 $Y2=2.44
r164 37 45 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.57 $Y=1.525
+ $X2=1.57 $Y2=1.392
r165 37 38 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.57 $Y=1.525
+ $X2=1.57 $Y2=2.32
r166 35 54 12.1487 $w=2.38e-07 $l=2.53e-07 $layer=LI1_cond $X=1.317 $Y=2.44
+ $X2=1.57 $Y2=2.44
r167 35 51 0.0960369 $w=2.38e-07 $l=2e-09 $layer=LI1_cond $X=1.317 $Y=2.44
+ $X2=1.315 $Y2=2.44
r168 31 45 11.7419 $w=2.63e-07 $l=2.7e-07 $layer=LI1_cond $X=1.3 $Y=1.392
+ $X2=1.57 $Y2=1.392
r169 31 33 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.3 $Y=1.26
+ $X2=1.3 $Y2=1.085
r170 29 30 41.3838 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=2.207 $Y=1.79
+ $X2=2.207 $Y2=1.885
r171 25 67 24.0971 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.995 $Y=1.885
+ $X2=3.995 $Y2=1.652
r172 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.995 $Y=1.885
+ $X2=3.995 $Y2=2.17
r173 24 66 24.0971 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.73 $Y=1.42
+ $X2=3.73 $Y2=1.652
r174 23 24 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=3.73 $Y=1.26
+ $X2=3.73 $Y2=1.42
r175 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.655 $Y=1.185
+ $X2=3.73 $Y2=1.26
r176 21 22 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.655 $Y=1.185
+ $X2=3.235 $Y2=1.185
r177 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.16 $Y=1.11
+ $X2=3.235 $Y2=1.185
r178 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.16 $Y=1.11
+ $X2=3.16 $Y2=0.715
r179 17 30 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.215 $Y=2.38
+ $X2=2.215 $Y2=1.885
r180 13 28 20.4101 $w=1.5e-07 $l=8.57321e-08 $layer=POLY_cond $X=2.2 $Y=1.41
+ $X2=2.177 $Y2=1.335
r181 13 29 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.2 $Y=1.41 $X2=2.2
+ $Y2=1.79
r182 9 28 20.4101 $w=1.5e-07 $l=8.52936e-08 $layer=POLY_cond $X=2.155 $Y=1.26
+ $X2=2.177 $Y2=1.335
r183 9 11 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.155 $Y=1.26
+ $X2=2.155 $Y2=0.74
r184 8 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.335
+ $X2=1.72 $Y2=1.335
r185 7 28 5.30422 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=2.08 $Y=1.335
+ $X2=2.177 $Y2=1.335
r186 7 8 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.08 $Y=1.335
+ $X2=1.885 $Y2=1.335
r187 2 51 300 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=2 $X=1.165
+ $Y=2.12 $X2=1.315 $Y2=2.405
r188 1 33 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.49 $X2=1.3 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%A_27_136# 1 2 8 9 11 14 19 24 25 28 29 31 33
+ 34
c82 34 0 1.4235e-19 $X=0.272 $Y=2.1
c83 28 0 8.07505e-20 $X=2.68 $Y=1.385
c84 24 0 1.8903e-19 $X=2.515 $Y=0.665
c85 14 0 2.97788e-19 $X=2.77 $Y=0.715
r86 33 34 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=2.265
+ $X2=0.272 $Y2=2.1
r87 31 34 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.185 $Y=1.25
+ $X2=0.185 $Y2=2.1
r88 29 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.385
+ $X2=2.68 $Y2=1.55
r89 29 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.385
+ $X2=2.68 $Y2=1.22
r90 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.385 $X2=2.68 $Y2=1.385
r91 26 28 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.68 $Y=0.75
+ $X2=2.68 $Y2=1.385
r92 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.515 $Y=0.665
+ $X2=2.68 $Y2=0.75
r93 24 25 135.048 $w=1.68e-07 $l=2.07e-06 $layer=LI1_cond $X=2.515 $Y=0.665
+ $X2=0.445 $Y2=0.665
r94 17 31 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=0.272 $Y=1.078
+ $X2=0.272 $Y2=1.25
r95 17 19 4.10871 $w=3.43e-07 $l=1.23e-07 $layer=LI1_cond $X=0.272 $Y=1.078
+ $X2=0.272 $Y2=0.955
r96 16 25 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.272 $Y=0.75
+ $X2=0.445 $Y2=0.665
r97 16 19 6.84785 $w=3.43e-07 $l=2.05e-07 $layer=LI1_cond $X=0.272 $Y=0.75
+ $X2=0.272 $Y2=0.955
r98 14 36 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.77 $Y=0.715
+ $X2=2.77 $Y2=1.22
r99 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.75 $Y=1.885
+ $X2=2.75 $Y2=2.46
r100 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.75 $Y=1.795 $X2=2.75
+ $Y2=1.885
r101 8 37 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=2.75 $Y=1.795
+ $X2=2.75 $Y2=1.55
r102 2 33 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r103 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%A_343_74# 1 2 7 9 12 14 15 21 24 25 29 31 32
+ 34 36 38
c107 31 0 6.57199e-20 $X=4.1 $Y=0.34
c108 24 0 1.29216e-19 $X=2.14 $Y=1.71
c109 15 0 1.68572e-19 $X=2.055 $Y=1.005
c110 12 0 1.87089e-19 $X=4.12 $Y=0.505
c111 7 0 8.07505e-20 $X=3.17 $Y=1.885
r112 36 39 4.98354 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.2 $Y=1.635
+ $X2=3.2 $Y2=1.795
r113 36 38 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=1.635
+ $X2=3.2 $Y2=1.47
r114 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.635 $X2=3.22 $Y2=1.635
r115 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.1
+ $Y=0.34 $X2=4.1 $Y2=0.34
r116 29 31 42.1794 $w=2.48e-07 $l=9.15e-07 $layer=LI1_cond $X=3.185 $Y=0.38
+ $X2=4.1 $Y2=0.38
r117 27 29 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.1 $Y=0.505
+ $X2=3.185 $Y2=0.38
r118 27 38 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=3.1 $Y=0.505
+ $X2=3.1 $Y2=1.47
r119 26 34 2.76166 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.225 $Y=1.795
+ $X2=2.025 $Y2=1.795
r120 25 39 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.015 $Y=1.795
+ $X2=3.2 $Y2=1.795
r121 25 26 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.015 $Y=1.795
+ $X2=2.225 $Y2=1.795
r122 24 34 3.70735 $w=2.5e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.14 $Y=1.71
+ $X2=2.025 $Y2=1.795
r123 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.14 $Y=1.09
+ $X2=2.14 $Y2=1.71
r124 19 34 3.70735 $w=2.5e-07 $l=1.00995e-07 $layer=LI1_cond $X=1.99 $Y=1.88
+ $X2=2.025 $Y2=1.795
r125 19 21 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.99 $Y=1.88
+ $X2=1.99 $Y2=2.12
r126 15 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.055 $Y=1.005
+ $X2=2.14 $Y2=1.09
r127 15 17 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.055 $Y=1.005
+ $X2=1.86 $Y2=1.005
r128 12 32 20.7597 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=4.12 $Y=0.505
+ $X2=4.155 $Y2=0.34
r129 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.12 $Y=0.505
+ $X2=4.12 $Y2=0.825
r130 7 37 52.2586 $w=2.99e-07 $l=2.73861e-07 $layer=POLY_cond $X=3.17 $Y=1.885
+ $X2=3.22 $Y2=1.635
r131 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.17 $Y=1.885
+ $X2=3.17 $Y2=2.46
r132 2 21 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.96 $X2=1.99 $Y2=2.12
r133 1 17 182 $w=1.7e-07 $l=7.03776e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.37 $X2=1.86 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%A_887_270# 1 2 7 9 12 16 18 20 23 25 27 30
+ 33 34 36 39 42 43 47 50 53 54 58 59 63 65 66 68 76
c155 58 0 1.78677e-19 $X=6.87 $Y=1.63
c156 43 0 3.16539e-20 $X=4.775 $Y=1.805
c157 12 0 6.57199e-20 $X=4.58 $Y=0.825
r158 73 74 12.6842 $w=3.61e-07 $l=9.5e-08 $layer=POLY_cond $X=6.555 $Y=1.532
+ $X2=6.65 $Y2=1.532
r159 72 73 47.3989 $w=3.61e-07 $l=3.55e-07 $layer=POLY_cond $X=6.2 $Y=1.532
+ $X2=6.555 $Y2=1.532
r160 71 72 10.0139 $w=3.61e-07 $l=7.5e-08 $layer=POLY_cond $X=6.125 $Y=1.532
+ $X2=6.2 $Y2=1.532
r161 69 76 46.0637 $w=3.61e-07 $l=3.45e-07 $layer=POLY_cond $X=6.79 $Y=1.532
+ $X2=7.135 $Y2=1.532
r162 69 74 18.6925 $w=3.61e-07 $l=1.4e-07 $layer=POLY_cond $X=6.79 $Y=1.532
+ $X2=6.65 $Y2=1.532
r163 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.79
+ $Y=1.465 $X2=6.79 $Y2=1.465
r164 61 63 5.3159 $w=4.93e-07 $l=2.2e-07 $layer=LI1_cond $X=5.35 $Y=0.597
+ $X2=5.57 $Y2=0.597
r165 58 68 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=1.63
+ $X2=6.87 $Y2=1.465
r166 58 59 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.87 $Y=1.63
+ $X2=6.87 $Y2=2.24
r167 55 66 4.59089 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.655 $Y=2.325
+ $X2=5.452 $Y2=2.325
r168 54 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.785 $Y=2.325
+ $X2=6.87 $Y2=2.24
r169 54 55 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=6.785 $Y=2.325
+ $X2=5.655 $Y2=2.325
r170 53 65 3.27229 $w=2.87e-07 $l=1.54771e-07 $layer=LI1_cond $X=5.57 $Y=1.72
+ $X2=5.452 $Y2=1.805
r171 52 63 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=5.57 $Y=0.845
+ $X2=5.57 $Y2=0.597
r172 52 53 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=5.57 $Y=0.845
+ $X2=5.57 $Y2=1.72
r173 48 66 2.39067 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.452 $Y=2.41
+ $X2=5.452 $Y2=2.325
r174 48 50 11.5244 $w=4.03e-07 $l=4.05e-07 $layer=LI1_cond $X=5.452 $Y=2.41
+ $X2=5.452 $Y2=2.815
r175 45 66 2.39067 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.452 $Y=2.24
+ $X2=5.452 $Y2=2.325
r176 45 47 7.25612 $w=4.03e-07 $l=2.55e-07 $layer=LI1_cond $X=5.452 $Y=2.24
+ $X2=5.452 $Y2=1.985
r177 44 65 3.27229 $w=2.87e-07 $l=8.5e-08 $layer=LI1_cond $X=5.452 $Y=1.89
+ $X2=5.452 $Y2=1.805
r178 44 47 2.70326 $w=4.03e-07 $l=9.5e-08 $layer=LI1_cond $X=5.452 $Y=1.89
+ $X2=5.452 $Y2=1.985
r179 42 65 3.2872 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=5.25 $Y=1.805
+ $X2=5.452 $Y2=1.805
r180 42 43 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.25 $Y=1.805
+ $X2=4.775 $Y2=1.805
r181 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.61
+ $Y=1.515 $X2=4.61 $Y2=1.515
r182 37 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.61 $Y=1.72
+ $X2=4.775 $Y2=1.805
r183 37 39 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.61 $Y=1.72
+ $X2=4.61 $Y2=1.515
r184 34 36 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.155 $Y=1.885
+ $X2=7.155 $Y2=2.46
r185 33 34 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.155 $Y=1.795
+ $X2=7.155 $Y2=1.885
r186 32 76 2.67036 $w=3.61e-07 $l=2e-08 $layer=POLY_cond $X=7.155 $Y=1.532
+ $X2=7.135 $Y2=1.532
r187 32 33 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.155 $Y=1.63
+ $X2=7.155 $Y2=1.795
r188 28 76 23.3725 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.135 $Y=1.3
+ $X2=7.135 $Y2=1.532
r189 28 30 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.135 $Y=1.3
+ $X2=7.135 $Y2=0.79
r190 25 74 23.3725 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.65 $Y=1.765
+ $X2=6.65 $Y2=1.532
r191 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.65 $Y=1.765
+ $X2=6.65 $Y2=2.4
r192 21 73 23.3725 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.555 $Y=1.3
+ $X2=6.555 $Y2=1.532
r193 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.555 $Y=1.3
+ $X2=6.555 $Y2=0.74
r194 18 72 23.3725 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.2 $Y=1.765
+ $X2=6.2 $Y2=1.532
r195 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.2 $Y=1.765
+ $X2=6.2 $Y2=2.4
r196 14 71 23.3725 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.125 $Y=1.3
+ $X2=6.125 $Y2=1.532
r197 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.125 $Y=1.3
+ $X2=6.125 $Y2=0.74
r198 10 40 38.7595 $w=2.78e-07 $l=1.77059e-07 $layer=POLY_cond $X=4.58 $Y=1.35
+ $X2=4.605 $Y2=1.515
r199 10 12 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.58 $Y=1.35
+ $X2=4.58 $Y2=0.825
r200 7 40 74.3026 $w=2.78e-07 $l=4.08044e-07 $layer=POLY_cond $X=4.525 $Y=1.885
+ $X2=4.605 $Y2=1.515
r201 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.525 $Y=1.885
+ $X2=4.525 $Y2=2.17
r202 2 50 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.84 $X2=5.415 $Y2=2.815
r203 2 47 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.84 $X2=5.415 $Y2=1.985
r204 1 61 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=5.21
+ $Y=0.37 $X2=5.35 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%A_647_79# 1 2 7 9 10 12 13 18 19 20 23 31
c80 10 0 1.15783e-19 $X=5.19 $Y=1.765
r81 29 31 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.64 $Y=2.135
+ $X2=3.77 $Y2=2.135
r82 26 28 7.64303 $w=4.23e-07 $l=2.65e-07 $layer=LI1_cond $X=3.64 $Y=0.955
+ $X2=3.905 $Y2=0.955
r83 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.15
+ $Y=1.385 $X2=5.15 $Y2=1.385
r84 21 23 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=5.15 $Y=1.185 $X2=5.15
+ $Y2=1.385
r85 20 28 9.26383 $w=4.23e-07 $l=2.26164e-07 $layer=LI1_cond $X=4.07 $Y=1.1
+ $X2=3.905 $Y2=0.955
r86 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.985 $Y=1.1
+ $X2=5.15 $Y2=1.185
r87 19 20 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=4.985 $Y=1.1
+ $X2=4.07 $Y2=1.1
r88 18 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=2.05
+ $X2=3.64 $Y2=2.135
r89 17 26 6.11956 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.64 $Y=1.185
+ $X2=3.64 $Y2=0.955
r90 17 18 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.64 $Y=1.185
+ $X2=3.64 $Y2=2.05
r91 13 29 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=2.135
+ $X2=3.64 $Y2=2.135
r92 13 15 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.555 $Y=2.135
+ $X2=3.395 $Y2=2.135
r93 10 24 77.2841 $w=2.7e-07 $l=3.995e-07 $layer=POLY_cond $X=5.19 $Y=1.765
+ $X2=5.15 $Y2=1.385
r94 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.19 $Y=1.765
+ $X2=5.19 $Y2=2.4
r95 7 24 38.9026 $w=2.7e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.135 $Y=1.22
+ $X2=5.15 $Y2=1.385
r96 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.135 $Y=1.22 $X2=5.135
+ $Y2=0.74
r97 2 31 600 $w=1.7e-07 $l=6.06218e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=1.96 $X2=3.77 $Y2=2.135
r98 2 15 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=1.96 $X2=3.395 $Y2=2.135
r99 1 28 91 $w=1.7e-07 $l=8.83487e-07 $layer=licon1_NDIFF $count=2 $X=3.235
+ $Y=0.395 $X2=3.905 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%A_1442_94# 1 2 7 9 12 14 16 19 21 24 28 31
+ 34 40 43 44
c64 34 0 1.28661e-19 $X=7.38 $Y=2.105
c65 24 0 1.83282e-19 $X=8.615 $Y=1.542
c66 21 0 1.78677e-19 $X=8.075 $Y=1.485
r67 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.99
+ $Y=1.485 $X2=7.99 $Y2=1.485
r68 38 44 1.17559 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.545 $Y=1.485
+ $X2=7.38 $Y2=1.485
r69 38 40 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.545 $Y=1.485
+ $X2=7.99 $Y2=1.485
r70 34 36 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.38 $Y=2.105
+ $X2=7.38 $Y2=2.815
r71 32 44 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=1.65
+ $X2=7.38 $Y2=1.485
r72 32 34 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=7.38 $Y=1.65
+ $X2=7.38 $Y2=2.105
r73 31 44 5.36902 $w=3.15e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.365 $Y=1.32
+ $X2=7.38 $Y2=1.485
r74 31 43 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=1.13
r75 26 43 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.35 $Y=0.965
+ $X2=7.35 $Y2=1.13
r76 26 28 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=7.35 $Y=0.965
+ $X2=7.35 $Y2=0.615
r77 24 25 1.22959 $w=3.92e-07 $l=1e-08 $layer=POLY_cond $X=8.615 $Y=1.542
+ $X2=8.625 $Y2=1.542
r78 23 24 51.6429 $w=3.92e-07 $l=4.2e-07 $layer=POLY_cond $X=8.195 $Y=1.542
+ $X2=8.615 $Y2=1.542
r79 22 23 3.68878 $w=3.92e-07 $l=3e-08 $layer=POLY_cond $X=8.165 $Y=1.542
+ $X2=8.195 $Y2=1.542
r80 21 41 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=8.075 $Y=1.485
+ $X2=7.99 $Y2=1.485
r81 21 22 12.4127 $w=3.92e-07 $l=1.15022e-07 $layer=POLY_cond $X=8.075 $Y=1.485
+ $X2=8.165 $Y2=1.542
r82 17 25 25.3688 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.625 $Y=1.32
+ $X2=8.625 $Y2=1.542
r83 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.625 $Y=1.32
+ $X2=8.625 $Y2=0.74
r84 14 24 25.3688 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=1.542
r85 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=2.4
r86 10 23 25.3688 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.195 $Y=1.32
+ $X2=8.195 $Y2=1.542
r87 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.195 $Y=1.32
+ $X2=8.195 $Y2=0.74
r88 7 22 25.3688 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=1.542
r89 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=2.4
r90 2 36 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.96 $X2=7.38 $Y2=2.815
r91 2 34 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.96 $X2=7.38 $Y2=2.105
r92 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.21
+ $Y=0.47 $X2=7.35 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%VPWR 1 2 3 4 5 6 7 26 30 34 40 44 48 52 54
+ 59 60 62 63 64 66 78 86 90 96 99 102 105 109
r98 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r99 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r100 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r101 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 94 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r104 94 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r106 91 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.9 $Y2=3.33
r107 91 93 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r108 90 108 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.937 $Y2=3.33
r109 90 93 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.4 $Y2=3.33
r110 89 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 86 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.9 $Y2=3.33
r113 86 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 85 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r116 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r117 82 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.14 $Y=3.33
+ $X2=6.015 $Y2=3.33
r118 82 84 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.14 $Y=3.33
+ $X2=6.48 $Y2=3.33
r119 81 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r120 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 78 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=6.015 $Y2=3.33
r122 78 80 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 74 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=2.525 $Y2=3.33
r124 74 76 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=2.69 $Y=3.33 $X2=4.56
+ $Y2=3.33
r125 73 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r126 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r127 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r128 70 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 69 72 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r130 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 67 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r132 67 69 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 66 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.525 $Y2=3.33
r134 66 72 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=3.33 $X2=2.16
+ $Y2=3.33
r135 64 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r136 64 100 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=2.64 $Y2=3.33
r137 64 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 62 84 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.48 $Y2=3.33
r139 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.875 $Y2=3.33
r140 61 88 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.04 $Y=3.33 $X2=7.44
+ $Y2=3.33
r141 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.04 $Y=3.33
+ $X2=6.875 $Y2=3.33
r142 59 76 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 59 60 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.875 $Y2=3.33
r144 58 80 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r145 58 60 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=5.08 $Y=3.33
+ $X2=4.875 $Y2=3.33
r146 54 57 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=2.815
r147 52 108 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.937 $Y2=3.33
r148 52 57 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.88 $Y2=2.815
r149 48 51 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.9 $Y=1.985
+ $X2=7.9 $Y2=2.815
r150 46 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=3.245
+ $X2=7.9 $Y2=3.33
r151 46 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.9 $Y=3.245 $X2=7.9
+ $Y2=2.815
r152 42 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=3.33
r153 42 44 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=2.78
r154 38 102 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=3.245
+ $X2=6.015 $Y2=3.33
r155 38 40 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=6.015 $Y=3.245
+ $X2=6.015 $Y2=2.78
r156 34 37 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=4.875 $Y=2.155
+ $X2=4.875 $Y2=2.495
r157 32 60 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=3.245
+ $X2=4.875 $Y2=3.33
r158 32 37 21.0813 $w=4.08e-07 $l=7.5e-07 $layer=LI1_cond $X=4.875 $Y=3.245
+ $X2=4.875 $Y2=2.495
r159 28 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=3.33
r160 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=2.815
r161 24 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r162 24 26 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.405
r163 7 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=2.815
r164 7 54 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=1.985
r165 6 51 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.94 $Y2=2.815
r166 6 48 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.94 $Y2=1.985
r167 5 44 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=6.725
+ $Y=1.84 $X2=6.875 $Y2=2.78
r168 4 40 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.975 $Y2=2.78
r169 3 37 300 $w=1.7e-07 $l=6.58293e-07 $layer=licon1_PDIFF $count=2 $X=4.6
+ $Y=1.96 $X2=4.875 $Y2=2.495
r170 3 34 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.96 $X2=4.875 $Y2=2.155
r171 2 30 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.96 $X2=2.525 $Y2=2.815
r172 1 26 300 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=2 $X=0.665
+ $Y=2.12 $X2=0.815 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%Q 1 2 7 9 13 20 23 24
r42 23 24 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6 $Y=1.295 $X2=6
+ $Y2=1.665
r43 22 24 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6 $Y=1.8 $X2=6
+ $Y2=1.665
r44 19 20 1.44055 $w=2.78e-07 $l=3.5e-08 $layer=LI1_cond $X=6.34 $Y=0.99
+ $X2=6.375 $Y2=0.99
r45 16 23 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=1.13 $X2=6
+ $Y2=1.295
r46 15 19 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=6 $Y=0.99 $X2=6.34
+ $Y2=0.99
r47 15 16 1.89134 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=6 $Y=0.99 $X2=6
+ $Y2=1.13
r48 11 20 1.16438 $w=2.6e-07 $l=1.4e-07 $layer=LI1_cond $X=6.375 $Y=0.85
+ $X2=6.375 $Y2=0.99
r49 11 13 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=6.375 $Y=0.85
+ $X2=6.375 $Y2=0.52
r50 7 22 6.87339 $w=2.7e-07 $l=1.83712e-07 $layer=LI1_cond $X=6.115 $Y=1.935
+ $X2=6 $Y2=1.8
r51 7 9 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.115 $Y=1.935
+ $X2=6.425 $Y2=1.935
r52 2 9 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.84 $X2=6.425 $Y2=1.985
r53 1 19 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=6.2
+ $Y=0.37 $X2=6.34 $Y2=0.95
r54 1 13 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=6.2
+ $Y=0.37 $X2=6.34 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%Q_N 1 2 9 13 14 15 16 24 33
r24 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.39 $Y=2.405
+ $X2=8.39 $Y2=2.775
r25 14 24 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=8.39 $Y=1.967
+ $X2=8.39 $Y2=1.985
r26 14 33 7.83357 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=8.39 $Y=1.967
+ $X2=8.39 $Y2=1.82
r27 14 15 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=8.39 $Y=2.052
+ $X2=8.39 $Y2=2.405
r28 14 24 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=8.39 $Y=2.052
+ $X2=8.39 $Y2=1.985
r29 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.41 $Y=1.13 $X2=8.41
+ $Y2=1.82
r30 7 13 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=8.37 $Y=1.005
+ $X2=8.37 $Y2=1.13
r31 7 9 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=8.37 $Y=1.005 $X2=8.37
+ $Y2=0.515
r32 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.24
+ $Y=1.84 $X2=8.39 $Y2=2.815
r33 2 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.24
+ $Y=1.84 $X2=8.39 $Y2=1.985
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.27
+ $Y=0.37 $X2=8.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_2%VGND 1 2 3 4 5 6 7 24 28 32 38 40 42 45 52
+ 53 55 56 58 59 60 62 86 90 97 103 107
c103 42 0 1.83282e-19 $X=8.84 $Y=0.515
c104 24 0 1.15783e-19 $X=4.82 $Y=0.76
r105 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r106 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r107 97 100 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0
+ $X2=0.79 $Y2=0.325
r108 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r109 94 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r110 94 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r111 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r112 91 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0
+ $X2=7.91 $Y2=0
r113 91 93 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=8.4
+ $Y2=0
r114 90 106 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.897 $Y2=0
r115 90 93 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=0 $X2=8.4
+ $Y2=0
r116 89 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r117 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r118 86 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.91 $Y2=0
r119 86 88 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r120 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r121 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r122 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r123 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r124 75 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r125 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r126 73 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r127 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r128 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r129 70 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r130 69 72 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r131 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r132 67 97 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r133 67 69 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r134 65 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r135 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r136 62 97 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r137 62 64 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r138 60 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r139 60 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=2.64 $Y2=0
r140 60 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r141 58 84 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.675 $Y=0
+ $X2=6.48 $Y2=0
r142 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.84
+ $Y2=0
r143 57 88 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.44 $Y2=0
r144 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0 $X2=6.84
+ $Y2=0
r145 55 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=5.52 $Y2=0
r146 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.825 $Y=0 $X2=5.95
+ $Y2=0
r147 54 84 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=6.48 $Y2=0
r148 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.075 $Y=0 $X2=5.95
+ $Y2=0
r149 52 78 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.63 $Y=0 $X2=4.56
+ $Y2=0
r150 52 53 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=4.63 $Y=0 $X2=4.822
+ $Y2=0
r151 51 81 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=5.015 $Y=0
+ $X2=5.52 $Y2=0
r152 51 53 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=5.015 $Y=0
+ $X2=4.822 $Y2=0
r153 45 72 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=0
+ $X2=2.16 $Y2=0
r154 45 49 10.5505 $w=3.53e-07 $l=3.25e-07 $layer=LI1_cond $X=2.462 $Y=0
+ $X2=2.462 $Y2=0.325
r155 45 75 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=2.462 $Y=0 $X2=2.64
+ $Y2=0
r156 40 106 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.897 $Y2=0
r157 40 42 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.84 $Y2=0.515
r158 36 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r159 36 38 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.515
r160 32 34 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.84 $Y=0.515
+ $X2=6.84 $Y2=0.965
r161 30 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0
r162 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0.515
r163 26 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0
r164 26 28 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0.515
r165 22 53 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.822 $Y=0.085
+ $X2=4.822 $Y2=0
r166 22 24 20.2052 $w=3.83e-07 $l=6.75e-07 $layer=LI1_cond $X=4.822 $Y=0.085
+ $X2=4.822 $Y2=0.76
r167 7 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r168 6 38 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.765
+ $Y=0.37 $X2=7.91 $Y2=0.515
r169 5 34 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=6.63
+ $Y=0.37 $X2=6.84 $Y2=0.965
r170 5 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.63
+ $Y=0.37 $X2=6.84 $Y2=0.515
r171 4 28 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=5.765
+ $Y=0.37 $X2=5.91 $Y2=0.515
r172 3 24 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.615 $X2=4.82 $Y2=0.76
r173 2 49 182 $w=1.7e-07 $l=2.51496e-07 $layer=licon1_NDIFF $count=1 $X=2.23
+ $Y=0.37 $X2=2.46 $Y2=0.325
r174 1 100 182 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.79 $Y2=0.325
.ends

