* File: sky130_fd_sc_hs__sedfxtp_1.pex.spice
* Created: Tue Sep  1 20:24:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%D 2 4 5 7 10 12 13 14 18 19
c44 18 0 4.24886e-20 $X=0.58 $Y=1.275
r45 18 20 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.275
+ $X2=0.575 $Y2=1.11
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.275 $X2=0.58 $Y2=1.275
r47 13 14 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.665
r48 13 19 0.606549 $w=3.78e-07 $l=2e-08 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.275
r49 10 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.64 $Y=0.58
+ $X2=0.64 $Y2=1.11
r50 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=2.245
+ $X2=0.495 $Y2=2.64
r51 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=2.155 $X2=0.495
+ $Y2=2.245
r52 4 12 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=0.495 $Y=2.155
+ $X2=0.495 $Y2=1.78
r53 2 12 41.5618 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=0.575 $Y=1.61
+ $X2=0.575 $Y2=1.78
r54 1 18 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.575 $Y=1.28
+ $X2=0.575 $Y2=1.275
r55 1 2 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=0.575 $Y=1.28 $X2=0.575
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_159_404# 1 2 7 9 12 14 20 21 22 23 24 25
+ 28 32 34 38 41 46
c116 41 0 9.40653e-20 $X=1.79 $Y=2.035
c117 23 0 4.24886e-20 $X=1.305 $Y=1.065
c118 21 0 1.72336e-19 $X=1.14 $Y=1.605
r119 39 46 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.22 $Y=1.685
+ $X2=2.45 $Y2=1.685
r120 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.685 $X2=2.22 $Y2=1.685
r121 36 38 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.22 $Y=1.95
+ $X2=2.22 $Y2=1.685
r122 35 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=2.035
+ $X2=1.79 $Y2=2.035
r123 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.055 $Y=2.035
+ $X2=2.22 $Y2=1.95
r124 34 35 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.055 $Y=2.035
+ $X2=1.875 $Y2=2.035
r125 30 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=2.12
+ $X2=1.79 $Y2=2.035
r126 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.79 $Y=2.12
+ $X2=1.79 $Y2=2.515
r127 26 28 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.765 $Y=0.98
+ $X2=1.765 $Y2=0.765
r128 24 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.035
+ $X2=1.79 $Y2=2.035
r129 24 25 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.705 $Y=2.035
+ $X2=1.305 $Y2=2.035
r130 22 26 14.8321 $w=1.01e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.64 $Y=1.065
+ $X2=1.765 $Y2=0.98
r131 22 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.64 $Y=1.065
+ $X2=1.305 $Y2=1.065
r132 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.605 $X2=1.14 $Y2=1.605
r133 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.95
+ $X2=1.305 $Y2=2.035
r134 18 20 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.14 $Y=1.95
+ $X2=1.14 $Y2=1.605
r135 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.15
+ $X2=1.305 $Y2=1.065
r136 17 20 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.14 $Y=1.15
+ $X2=1.14 $Y2=1.605
r137 16 21 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=1.14 $Y=2.02
+ $X2=1.14 $Y2=1.605
r138 14 16 79.2968 $w=1.55e-07 $l=3.05917e-07 $layer=POLY_cond $X=0.885 $Y=2.132
+ $X2=1.14 $Y2=2.02
r139 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=1.52
+ $X2=2.45 $Y2=1.685
r140 10 12 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.45 $Y=1.52
+ $X2=2.45 $Y2=0.765
r141 7 14 3.61756 $w=1.5e-07 $l=1.13e-07 $layer=POLY_cond $X=0.885 $Y=2.245
+ $X2=0.885 $Y2=2.132
r142 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.885 $Y=2.245
+ $X2=0.885 $Y2=2.64
r143 2 32 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=2.315 $X2=1.79 $Y2=2.515
r144 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.555 $X2=1.805 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%DE 3 5 6 10 11 13 14 16 17 18 19 21 23 28
+ 31 32 33
c90 33 0 9.40653e-20 $X=1.68 $Y=1.65
c91 32 0 1.3237e-19 $X=1.68 $Y=1.485
r92 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.485
+ $X2=1.68 $Y2=1.65
r93 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.485 $X2=1.68 $Y2=1.485
r94 28 32 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.485
r95 25 27 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=1.74 $Y=2.165
+ $X2=2.015 $Y2=2.165
r96 19 21 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.695 $Y=2.24
+ $X2=2.695 $Y2=2.635
r97 18 27 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.09 $Y=2.165
+ $X2=2.015 $Y2=2.165
r98 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.62 $Y=2.165
+ $X2=2.695 $Y2=2.24
r99 17 18 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.62 $Y=2.165
+ $X2=2.09 $Y2=2.165
r100 14 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.02 $Y=1.05
+ $X2=2.02 $Y2=1.125
r101 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.02 $Y=1.05
+ $X2=2.02 $Y2=0.765
r102 11 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.015 $Y=2.24
+ $X2=2.015 $Y2=2.165
r103 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.015 $Y=2.24
+ $X2=2.015 $Y2=2.635
r104 10 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.74 $Y=2.09
+ $X2=1.74 $Y2=2.165
r105 10 33 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.74 $Y=2.09
+ $X2=1.74 $Y2=1.65
r106 7 23 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.68 $Y=1.125
+ $X2=2.02 $Y2=1.125
r107 7 31 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.68 $Y=1.2
+ $X2=1.68 $Y2=1.485
r108 5 7 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.125
+ $X2=1.68 $Y2=1.125
r109 5 6 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.515 $Y=1.125
+ $X2=1.105 $Y2=1.125
r110 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.03 $Y=1.05
+ $X2=1.105 $Y2=1.125
r111 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.03 $Y=1.05 $X2=1.03
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_547_301# 1 2 9 12 13 15 16 18 19 20 21
+ 23 25 26 33 36 40 43 44 45 51 52 58 59 67
c238 52 0 8.71884e-20 $X=14.16 $Y=1.665
c239 44 0 7.68314e-20 $X=14.015 $Y=1.665
c240 13 0 1.85697e-19 $X=3.085 $Y=2.24
r241 57 59 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.9 $Y=1.67
+ $X2=3.085 $Y2=1.67
r242 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.9
+ $Y=1.67 $X2=2.9 $Y2=1.67
r243 54 57 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.84 $Y=1.67 $X2=2.9
+ $Y2=1.67
r244 52 67 6.51792 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=14.165 $Y=1.665
+ $X2=14.165 $Y2=1.55
r245 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=1.665
+ $X2=14.16 $Y2=1.665
r246 48 58 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.64 $Y=1.67
+ $X2=2.9 $Y2=1.67
r247 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r248 45 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r249 44 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.015 $Y=1.665
+ $X2=14.16 $Y2=1.665
r250 44 45 13.8985 $w=1.4e-07 $l=1.123e-05 $layer=MET1_cond $X=14.015 $Y=1.665
+ $X2=2.785 $Y2=1.665
r251 42 67 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=14.2 $Y=0.81
+ $X2=14.2 $Y2=1.55
r252 40 42 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=14.105 $Y=0.58
+ $X2=14.105 $Y2=0.81
r253 36 43 5.46396 $w=2.85e-07 $l=1.73043e-07 $layer=LI1_cond $X=14.165 $Y=2.075
+ $X2=14.12 $Y2=2.227
r254 35 52 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=14.165 $Y=1.67
+ $X2=14.165 $Y2=1.665
r255 35 36 19.4475 $w=2.38e-07 $l=4.05e-07 $layer=LI1_cond $X=14.165 $Y=1.67
+ $X2=14.165 $Y2=2.075
r256 31 43 5.46396 $w=2.85e-07 $l=1.53e-07 $layer=LI1_cond $X=14.12 $Y=2.38
+ $X2=14.12 $Y2=2.227
r257 31 33 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=14.12 $Y=2.38
+ $X2=14.12 $Y2=2.465
r258 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.23
+ $Y=2.215 $X2=13.23 $Y2=2.215
r259 26 43 1.09951 $w=3.05e-07 $l=1.65e-07 $layer=LI1_cond $X=13.955 $Y=2.227
+ $X2=14.12 $Y2=2.227
r260 26 28 27.3941 $w=3.03e-07 $l=7.25e-07 $layer=LI1_cond $X=13.955 $Y=2.227
+ $X2=13.23 $Y2=2.227
r261 25 29 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=13.29 $Y=2.05
+ $X2=13.23 $Y2=2.215
r262 24 25 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=13.29 $Y=1.015
+ $X2=13.29 $Y2=2.05
r263 21 29 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=13.185 $Y=2.465
+ $X2=13.23 $Y2=2.215
r264 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.185 $Y=2.465
+ $X2=13.185 $Y2=2.75
r265 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.215 $Y=0.94
+ $X2=13.29 $Y2=1.015
r266 19 20 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=13.215 $Y=0.94
+ $X2=12.825 $Y2=0.94
r267 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.75 $Y=0.865
+ $X2=12.825 $Y2=0.94
r268 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.75 $Y=0.865
+ $X2=12.75 $Y2=0.58
r269 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.085 $Y=2.24
+ $X2=3.085 $Y2=2.635
r270 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.085 $Y=2.15
+ $X2=3.085 $Y2=2.24
r271 11 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.835
+ $X2=3.085 $Y2=1.67
r272 11 12 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=3.085 $Y=1.835
+ $X2=3.085 $Y2=2.15
r273 7 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.505
+ $X2=2.84 $Y2=1.67
r274 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.84 $Y=1.505
+ $X2=2.84 $Y2=0.765
r275 2 33 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=13.97
+ $Y=2.32 $X2=14.12 $Y2=2.465
r276 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.95
+ $Y=0.37 $X2=14.09 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_639_85# 1 2 7 9 10 11 12 14 17 18 21 22
+ 27 28 30 31 35 36 41 43 47
c114 41 0 1.30585e-19 $X=4.41 $Y=0.805
c115 36 0 1.64952e-19 $X=5.655 $Y=1.58
r116 44 47 4.60989 $w=4.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.1 $Y=2.495
+ $X2=4.285 $Y2=2.495
r117 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.655
+ $Y=1.58 $X2=5.655 $Y2=1.58
r118 33 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.655 $Y=1.915
+ $X2=5.655 $Y2=1.58
r119 32 43 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.185 $Y=2 $X2=4.045
+ $Y2=2
r120 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.49 $Y=2
+ $X2=5.655 $Y2=1.915
r121 31 32 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=5.49 $Y=2
+ $X2=4.185 $Y2=2
r122 30 44 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=4.1 $Y=2.255 $X2=4.1
+ $Y2=2.495
r123 29 43 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=4.1 $Y=2.085
+ $X2=4.045 $Y2=2
r124 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.1 $Y=2.085
+ $X2=4.1 $Y2=2.255
r125 27 28 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.995
+ $Y=1.78 $X2=3.995 $Y2=1.78
r126 25 43 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=1.915
+ $X2=4.045 $Y2=2
r127 25 27 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=4.045 $Y=1.915
+ $X2=4.045 $Y2=1.78
r128 24 27 31.6922 $w=2.78e-07 $l=7.7e-07 $layer=LI1_cond $X=4.045 $Y=1.01
+ $X2=4.045 $Y2=1.78
r129 21 22 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.995
+ $Y=0.42 $X2=3.995 $Y2=0.42
r130 19 41 10.3862 $w=4.03e-07 $l=3.65e-07 $layer=LI1_cond $X=4.045 $Y=0.807
+ $X2=4.41 $Y2=0.807
r131 19 24 2.89865 $w=2.8e-07 $l=2.03e-07 $layer=LI1_cond $X=4.045 $Y=0.807
+ $X2=4.045 $Y2=1.01
r132 19 21 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.045 $Y=0.605
+ $X2=4.045 $Y2=0.42
r133 18 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.655 $Y=1.92
+ $X2=5.655 $Y2=1.58
r134 16 28 101.42 $w=3.3e-07 $l=5.8e-07 $layer=POLY_cond $X=3.995 $Y=1.2
+ $X2=3.995 $Y2=1.78
r135 16 17 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.995 $Y=1.2
+ $X2=3.995 $Y2=1.125
r136 15 22 110.163 $w=3.3e-07 $l=6.3e-07 $layer=POLY_cond $X=3.995 $Y=1.05
+ $X2=3.995 $Y2=0.42
r137 15 17 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.995 $Y=1.05
+ $X2=3.995 $Y2=1.125
r138 12 18 50.3582 $w=2.68e-07 $l=3.15278e-07 $layer=POLY_cond $X=5.58 $Y=2.2
+ $X2=5.655 $Y2=1.92
r139 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.58 $Y=2.2
+ $X2=5.58 $Y2=2.595
r140 10 17 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.125
+ $X2=3.995 $Y2=1.125
r141 10 11 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.83 $Y=1.125
+ $X2=3.345 $Y2=1.125
r142 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.27 $Y=1.05
+ $X2=3.345 $Y2=1.125
r143 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.27 $Y=1.05 $X2=3.27
+ $Y2=0.765
r144 2 47 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=4.155
+ $Y=2.275 $X2=4.285 $Y2=2.495
r145 1 41 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.625 $X2=4.41 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%SCD 3 6 7 9 10 13
c46 13 0 1.14523e-19 $X=5.115 $Y=1.58
c47 3 0 1.30585e-19 $X=5.055 $Y=0.835
r48 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.58
+ $X2=5.115 $Y2=1.745
r49 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.58
+ $X2=5.115 $Y2=1.415
r50 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.58 $X2=5.115 $Y2=1.58
r51 10 14 9.25201 $w=3.53e-07 $l=2.85e-07 $layer=LI1_cond $X=5.102 $Y=1.295
+ $X2=5.102 $Y2=1.58
r52 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.19 $Y=2.2 $X2=5.19
+ $Y2=2.595
r53 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.19 $Y=2.11 $X2=5.19
+ $Y2=2.2
r54 6 16 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=5.19 $Y=2.11
+ $X2=5.19 $Y2=1.745
r55 3 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.055 $Y=0.835
+ $X2=5.055 $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%SCE 1 3 4 5 7 8 11 15 16 17 20 22 25
c86 25 0 5.07631e-20 $X=4.565 $Y=1.345
c87 22 0 1.14523e-19 $X=4.56 $Y=1.295
r88 25 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.345
+ $X2=4.565 $Y2=1.51
r89 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.345
+ $X2=4.565 $Y2=1.18
r90 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.565
+ $Y=1.345 $X2=4.565 $Y2=1.345
r91 18 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.415 $Y=0.255
+ $X2=5.415 $Y2=0.835
r92 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.34 $Y=0.18
+ $X2=5.415 $Y2=0.255
r93 16 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.34 $Y=0.18 $X2=4.7
+ $Y2=0.18
r94 15 27 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.625 $Y=0.835
+ $X2=4.625 $Y2=1.18
r95 12 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.625 $Y=0.255
+ $X2=4.7 $Y2=0.18
r96 12 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.625 $Y=0.255
+ $X2=4.625 $Y2=0.835
r97 9 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.51 $Y=2.99
+ $X2=4.51 $Y2=2.595
r98 8 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.51 $Y=2.2 $X2=4.51
+ $Y2=2.595
r99 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.51 $Y=2.11 $X2=4.51
+ $Y2=2.2
r100 7 28 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.51 $Y=2.11 $X2=4.51
+ $Y2=1.51
r101 4 9 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=4.42 $Y=3.105
+ $X2=4.51 $Y2=2.99
r102 4 5 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.42 $Y=3.105 $X2=3.61
+ $Y2=3.105
r103 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.535 $Y=3.03
+ $X2=3.61 $Y2=3.105
r104 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.535 $Y=3.03
+ $X2=3.535 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%CLK 1 3 4 6 7
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.495
+ $Y=1.385 $X2=6.495 $Y2=1.385
r34 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.495 $Y=1.295
+ $X2=6.495 $Y2=1.385
r35 4 10 64.88 $w=2.85e-07 $l=3.47793e-07 $layer=POLY_cond $X=6.55 $Y=1.705
+ $X2=6.492 $Y2=1.385
r36 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.55 $Y=1.705
+ $X2=6.55 $Y2=2.34
r37 1 10 38.666 $w=2.85e-07 $l=2.05925e-07 $layer=POLY_cond $X=6.4 $Y=1.22
+ $X2=6.492 $Y2=1.385
r38 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.4 $Y=1.22 $X2=6.4
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1492_74# 1 2 7 9 10 12 15 18 19 21 24 26
+ 27 28 33 34 37 40 41 43 46 47 48 50 51 52 53 55 56 58 60 64 65 68 72
c233 72 0 2.60684e-20 $X=12.84 $Y=1.39
c234 64 0 6.63657e-20 $X=8.575 $Y=2.17
c235 56 0 6.25838e-20 $X=11.76 $Y=1.635
c236 37 0 1.94394e-19 $X=9.17 $Y=0.85
c237 33 0 1.24564e-19 $X=8.49 $Y=1.82
c238 19 0 1.20815e-19 $X=12.765 $Y=2.465
r239 72 85 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.84 $Y=1.39
+ $X2=12.84 $Y2=1.555
r240 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.84
+ $Y=1.39 $X2=12.84 $Y2=1.39
r241 68 71 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=12.84 $Y=1.195
+ $X2=12.84 $Y2=1.39
r242 66 67 14.0135 $w=2.22e-07 $l=2.55e-07 $layer=LI1_cond $X=11.71 $Y=0.94
+ $X2=11.71 $Y2=1.195
r243 64 75 48.3612 $w=2.99e-07 $l=3e-07 $layer=POLY_cond $X=8.575 $Y=2.235
+ $X2=8.875 $Y2=2.235
r244 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.575
+ $Y=2.17 $X2=8.575 $Y2=2.17
r245 59 67 2.3025 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=11.86 $Y=1.195
+ $X2=11.71 $Y2=1.195
r246 58 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.675 $Y=1.195
+ $X2=12.84 $Y2=1.195
r247 58 59 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=12.675 $Y=1.195
+ $X2=11.86 $Y2=1.195
r248 56 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.76 $Y=1.635
+ $X2=11.76 $Y2=1.47
r249 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.76
+ $Y=1.635 $X2=11.76 $Y2=1.635
r250 53 67 4.30642 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.71 $Y=1.28
+ $X2=11.71 $Y2=1.195
r251 53 55 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=11.71 $Y=1.28
+ $X2=11.71 $Y2=1.635
r252 51 66 2.3025 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=11.56 $Y=0.94
+ $X2=11.71 $Y2=0.94
r253 51 52 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=11.56 $Y=0.94
+ $X2=11.02 $Y2=0.94
r254 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.935 $Y=0.855
+ $X2=11.02 $Y2=0.94
r255 49 50 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.935 $Y=0.425
+ $X2=10.935 $Y2=0.855
r256 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.85 $Y=0.34
+ $X2=10.935 $Y2=0.425
r257 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.85 $Y=0.34
+ $X2=10.34 $Y2=0.34
r258 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.255 $Y=0.425
+ $X2=10.34 $Y2=0.34
r259 45 46 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.255 $Y=0.425
+ $X2=10.255 $Y2=0.85
r260 44 65 2.15711 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.34 $Y=0.935
+ $X2=9.212 $Y2=0.935
r261 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.17 $Y=0.935
+ $X2=10.255 $Y2=0.85
r262 43 44 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=10.17 $Y=0.935
+ $X2=9.34 $Y2=0.935
r263 41 76 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=9.175 $Y=1.18
+ $X2=9.045 $Y2=1.18
r264 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.175
+ $Y=1.18 $X2=9.175 $Y2=1.18
r265 38 65 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=9.212 $Y=1.02
+ $X2=9.212 $Y2=0.935
r266 38 40 7.23101 $w=2.53e-07 $l=1.6e-07 $layer=LI1_cond $X=9.212 $Y=1.02
+ $X2=9.212 $Y2=1.18
r267 37 65 4.27425 $w=2.12e-07 $l=1.03899e-07 $layer=LI1_cond $X=9.17 $Y=0.85
+ $X2=9.212 $Y2=0.935
r268 36 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.17 $Y=0.425
+ $X2=9.17 $Y2=0.85
r269 35 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.575 $Y=0.34
+ $X2=8.49 $Y2=0.34
r270 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.085 $Y=0.34
+ $X2=9.17 $Y2=0.425
r271 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.085 $Y=0.34
+ $X2=8.575 $Y2=0.34
r272 32 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.49 $Y=0.425
+ $X2=8.49 $Y2=0.34
r273 32 33 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.49 $Y=0.425
+ $X2=8.49 $Y2=1.82
r274 28 63 9.54783 $w=2.3e-07 $l=1.8e-07 $layer=LI1_cond $X=8.535 $Y=1.99
+ $X2=8.535 $Y2=2.17
r275 28 33 9.87245 $w=2.3e-07 $l=1.91181e-07 $layer=LI1_cond $X=8.535 $Y=1.99
+ $X2=8.49 $Y2=1.82
r276 28 30 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=8.405 $Y=1.99
+ $X2=8.125 $Y2=1.99
r277 26 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=0.34
+ $X2=8.49 $Y2=0.34
r278 26 27 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.405 $Y=0.34
+ $X2=7.765 $Y2=0.34
r279 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.64 $Y=0.425
+ $X2=7.765 $Y2=0.34
r280 22 24 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.64 $Y=0.425
+ $X2=7.64 $Y2=0.515
r281 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.765 $Y=2.465
+ $X2=12.765 $Y2=2.75
r282 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.765 $Y=2.375
+ $X2=12.765 $Y2=2.465
r283 18 85 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=12.765 $Y=2.375
+ $X2=12.765 $Y2=1.555
r284 15 81 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=11.85 $Y=0.69
+ $X2=11.85 $Y2=1.47
r285 10 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.045 $Y=1.015
+ $X2=9.045 $Y2=1.18
r286 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.045 $Y=1.015
+ $X2=9.045 $Y2=0.695
r287 7 75 18.89 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=8.875 $Y=2.465
+ $X2=8.875 $Y2=2.235
r288 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.875 $Y=2.465
+ $X2=8.875 $Y2=2.75
r289 2 30 600 $w=1.7e-07 $l=2.12132e-07 $layer=licon1_PDIFF $count=1 $X=7.975
+ $Y=1.84 $X2=8.125 $Y2=1.99
r290 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.46
+ $Y=0.37 $X2=7.6 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1295_74# 1 2 9 11 13 15 16 20 22 25 26
+ 28 29 31 34 37 38 39 42 45 48 49 51 57 58 59 61 64 70 74
c200 58 0 1.20815e-19 $X=12.03 $Y=2.475
c201 57 0 2.75377e-20 $X=9.57 $Y=2.39
c202 51 0 3.8828e-20 $X=9.485 $Y=2.09
c203 26 0 7.11901e-20 $X=9.375 $Y=2.465
c204 25 0 1.24564e-19 $X=9.25 $Y=1.925
c205 20 0 1.94394e-19 $X=8.365 $Y=0.695
r206 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.3
+ $Y=1.59 $X2=12.3 $Y2=1.59
r207 71 74 7.48077 $w=2.83e-07 $l=1.85e-07 $layer=LI1_cond $X=12.115 $Y=1.592
+ $X2=12.3 $Y2=1.592
r208 69 70 2.83598 $w=3.98e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=1.96 $X2=7
+ $Y2=1.96
r209 67 69 4.03355 $w=3.98e-07 $l=1.4e-07 $layer=LI1_cond $X=6.775 $Y=1.96
+ $X2=6.915 $Y2=1.96
r210 60 71 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=12.115 $Y=1.735
+ $X2=12.115 $Y2=1.592
r211 60 61 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=12.115 $Y=1.735
+ $X2=12.115 $Y2=2.39
r212 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.03 $Y=2.475
+ $X2=12.115 $Y2=2.39
r213 58 59 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=12.03 $Y=2.475
+ $X2=9.655 $Y2=2.475
r214 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.57 $Y=2.39
+ $X2=9.655 $Y2=2.475
r215 56 57 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.57 $Y=2.22
+ $X2=9.57 $Y2=2.39
r216 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.34
+ $Y=2.09 $X2=9.34 $Y2=2.09
r217 51 56 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.485 $Y=2.09
+ $X2=9.57 $Y2=2.22
r218 51 53 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=9.485 $Y=2.09
+ $X2=9.34 $Y2=2.09
r219 48 70 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=7.225 $Y=1.995
+ $X2=7 $Y2=1.995
r220 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.225
+ $Y=1.995 $X2=7.225 $Y2=1.995
r221 45 69 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.915 $Y=1.76
+ $X2=6.915 $Y2=1.96
r222 44 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=1.01
+ $X2=6.915 $Y2=0.925
r223 44 45 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.915 $Y=1.01
+ $X2=6.915 $Y2=1.76
r224 40 64 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.615 $Y=0.925
+ $X2=6.915 $Y2=0.925
r225 40 42 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.615 $Y=0.84
+ $X2=6.615 $Y2=0.515
r226 36 49 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=7.225 $Y=1.765
+ $X2=7.225 $Y2=1.995
r227 36 37 13.5877 $w=2.4e-07 $l=9.08295e-08 $layer=POLY_cond $X=7.225 $Y=1.765
+ $X2=7.26 $Y2=1.69
r228 32 75 38.6443 $w=2.87e-07 $l=1.92678e-07 $layer=POLY_cond $X=12.36 $Y=1.425
+ $X2=12.3 $Y2=1.59
r229 32 34 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=12.36 $Y=1.425
+ $X2=12.36 $Y2=0.58
r230 29 75 60.4771 $w=2.87e-07 $l=3.28139e-07 $layer=POLY_cond $X=12.23 $Y=1.885
+ $X2=12.3 $Y2=1.59
r231 29 31 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.23 $Y=1.885
+ $X2=12.23 $Y2=2.46
r232 26 54 76.233 $w=2.71e-07 $l=3.9211e-07 $layer=POLY_cond $X=9.375 $Y=2.465
+ $X2=9.34 $Y2=2.09
r233 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.375 $Y=2.465
+ $X2=9.375 $Y2=2.75
r234 25 54 38.8824 $w=2.71e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.25 $Y=1.925
+ $X2=9.34 $Y2=2.09
r235 24 25 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=9.25 $Y=1.765
+ $X2=9.25 $Y2=1.925
r236 23 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.44 $Y=1.69
+ $X2=8.365 $Y2=1.69
r237 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.175 $Y=1.69
+ $X2=9.25 $Y2=1.765
r238 22 23 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=9.175 $Y=1.69
+ $X2=8.44 $Y2=1.69
r239 18 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.365 $Y=1.615
+ $X2=8.365 $Y2=1.69
r240 18 20 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=8.365 $Y=1.615
+ $X2=8.365 $Y2=0.695
r241 17 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.975 $Y=1.69
+ $X2=7.9 $Y2=1.69
r242 16 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.29 $Y=1.69
+ $X2=8.365 $Y2=1.69
r243 16 17 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=8.29 $Y=1.69
+ $X2=7.975 $Y2=1.69
r244 13 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.9 $Y=1.765
+ $X2=7.9 $Y2=1.69
r245 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.9 $Y=1.765
+ $X2=7.9 $Y2=2.4
r246 12 37 12.1617 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.46 $Y=1.69 $X2=7.26
+ $Y2=1.69
r247 11 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.825 $Y=1.69
+ $X2=7.9 $Y2=1.69
r248 11 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=7.825 $Y=1.69
+ $X2=7.46 $Y2=1.69
r249 7 37 13.5877 $w=2.4e-07 $l=1.58114e-07 $layer=POLY_cond $X=7.385 $Y=1.615
+ $X2=7.26 $Y2=1.69
r250 7 9 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=7.385 $Y=1.615
+ $X2=7.385 $Y2=0.74
r251 2 67 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.78 $X2=6.775 $Y2=1.96
r252 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.475
+ $Y=0.37 $X2=6.615 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1910_71# 1 2 9 12 13 15 19 20 22 23 25
+ 26 30 33 34 36 37 43 47 54 57
c113 36 0 6.25838e-20 $X=11.22 $Y=1.36
r114 49 50 5.82061 $w=2.62e-07 $l=1.25e-07 $layer=LI1_cond $X=10.595 $Y=1.36
+ $X2=10.72 $Y2=1.36
r115 45 47 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=10.55 $Y=2.095
+ $X2=10.72 $Y2=2.095
r116 41 54 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.73 $Y=1.32
+ $X2=9.805 $Y2=1.32
r117 41 51 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=9.73 $Y=1.32
+ $X2=9.625 $Y2=1.32
r118 40 43 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.73 $Y=1.32
+ $X2=9.895 $Y2=1.32
r119 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.73
+ $Y=1.32 $X2=9.73 $Y2=1.32
r120 37 57 12.8191 $w=2.82e-07 $l=7.5e-08 $layer=POLY_cond $X=11.22 $Y=1.317
+ $X2=11.295 $Y2=1.317
r121 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.22
+ $Y=1.36 $X2=11.22 $Y2=1.36
r122 34 50 3.69502 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.805 $Y=1.36
+ $X2=10.72 $Y2=1.36
r123 34 36 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=10.805 $Y=1.36
+ $X2=11.22 $Y2=1.36
r124 33 47 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.72 $Y=1.97
+ $X2=10.72 $Y2=2.095
r125 32 50 3.26844 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.72 $Y=1.525
+ $X2=10.72 $Y2=1.36
r126 32 33 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=10.72 $Y=1.525
+ $X2=10.72 $Y2=1.97
r127 28 49 3.26844 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.595 $Y=1.195
+ $X2=10.595 $Y2=1.36
r128 28 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.595 $Y=1.195
+ $X2=10.595 $Y2=0.81
r129 26 49 5.45986 $w=2.62e-07 $l=1.18427e-07 $layer=LI1_cond $X=10.51 $Y=1.28
+ $X2=10.595 $Y2=1.36
r130 26 43 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=10.51 $Y=1.28
+ $X2=9.895 $Y2=1.28
r131 23 57 33.3298 $w=2.82e-07 $l=2.88468e-07 $layer=POLY_cond $X=11.49 $Y=1.11
+ $X2=11.295 $Y2=1.317
r132 23 25 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=11.49 $Y=1.11
+ $X2=11.49 $Y2=0.69
r133 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.295 $Y=1.885
+ $X2=11.295 $Y2=2.46
r134 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.295 $Y=1.795
+ $X2=11.295 $Y2=1.885
r135 18 57 13.2911 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.295 $Y=1.525
+ $X2=11.295 $Y2=1.317
r136 18 19 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=11.295 $Y=1.525
+ $X2=11.295 $Y2=1.795
r137 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.805 $Y=2.465
+ $X2=9.805 $Y2=2.75
r138 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.805 $Y=2.375
+ $X2=9.805 $Y2=2.465
r139 11 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.805 $Y=1.485
+ $X2=9.805 $Y2=1.32
r140 11 12 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=9.805 $Y=1.485
+ $X2=9.805 $Y2=2.375
r141 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.625 $Y=1.155
+ $X2=9.625 $Y2=1.32
r142 7 9 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=9.625 $Y=1.155
+ $X2=9.625 $Y2=0.695
r143 2 45 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.4
+ $Y=1.99 $X2=10.55 $Y2=2.135
r144 1 30 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=10.455
+ $Y=0.37 $X2=10.595 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1688_97# 1 2 7 9 12 16 22 26 27 28 30 32
r98 30 32 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.3 $Y=1.665
+ $X2=10.135 $Y2=1.665
r99 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.3
+ $Y=1.665 $X2=10.3 $Y2=1.665
r100 27 28 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.075 $Y=2.39
+ $X2=9.075 $Y2=2.56
r101 25 26 1.34256 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.005 $Y=1.705
+ $X2=8.875 $Y2=1.705
r102 25 32 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=9.005 $Y=1.705
+ $X2=10.135 $Y2=1.705
r103 22 28 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.15 $Y=2.75
+ $X2=9.15 $Y2=2.56
r104 18 26 5.16603 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=8.92 $Y=1.79
+ $X2=8.875 $Y2=1.705
r105 18 27 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.92 $Y=1.79 $X2=8.92
+ $Y2=2.39
r106 14 26 5.16603 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=8.83 $Y=1.62
+ $X2=8.875 $Y2=1.705
r107 14 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=8.83 $Y=1.62
+ $X2=8.83 $Y2=0.76
r108 10 31 38.5562 $w=2.99e-07 $l=2.0106e-07 $layer=POLY_cond $X=10.38 $Y=1.5
+ $X2=10.3 $Y2=1.665
r109 10 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.38 $Y=1.5
+ $X2=10.38 $Y2=0.69
r110 7 31 52.2586 $w=2.99e-07 $l=2.62202e-07 $layer=POLY_cond $X=10.325 $Y=1.915
+ $X2=10.3 $Y2=1.665
r111 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.325 $Y=1.915
+ $X2=10.325 $Y2=2.41
r112 2 22 600 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_PDIFF $count=1 $X=8.95
+ $Y=2.54 $X2=9.15 $Y2=2.75
r113 1 16 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=8.44
+ $Y=0.485 $X2=8.83 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_2385_74# 1 2 9 12 13 15 16 17 18 20 21
+ 23 24 25 27 29 31 33 35 38 39 42 48 50
c144 25 0 1.37761e-19 $X=12.065 $Y=0.77
r145 55 56 2.23148 $w=4.32e-07 $l=2e-08 $layer=POLY_cond $X=13.875 $Y=1.335
+ $X2=13.895 $Y2=1.335
r146 51 55 10.5995 $w=4.32e-07 $l=9.5e-08 $layer=POLY_cond $X=13.78 $Y=1.335
+ $X2=13.875 $Y2=1.335
r147 50 53 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.78 $Y=1.215
+ $X2=13.78 $Y2=1.38
r148 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.78
+ $Y=1.215 $X2=13.78 $Y2=1.215
r149 42 53 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.7 $Y=1.735
+ $X2=13.7 $Y2=1.38
r150 40 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.345 $Y=1.82
+ $X2=13.26 $Y2=1.82
r151 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.615 $Y=1.82
+ $X2=13.7 $Y2=1.735
r152 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=13.615 $Y=1.82
+ $X2=13.345 $Y2=1.82
r153 38 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.26 $Y=1.735
+ $X2=13.26 $Y2=1.82
r154 37 38 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=13.26 $Y=0.94
+ $X2=13.26 $Y2=1.735
r155 36 47 11.3627 $w=3.06e-07 $l=3.78622e-07 $layer=LI1_cond $X=12.805 $Y=1.82
+ $X2=12.587 $Y2=2.105
r156 35 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.175 $Y=1.82
+ $X2=13.26 $Y2=1.82
r157 35 36 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.175 $Y=1.82
+ $X2=12.805 $Y2=1.82
r158 31 47 2.54614 $w=4.35e-07 $l=5.2e-08 $layer=LI1_cond $X=12.587 $Y=2.157
+ $X2=12.587 $Y2=2.105
r159 31 33 17.4324 $w=4.33e-07 $l=6.58e-07 $layer=LI1_cond $X=12.587 $Y=2.157
+ $X2=12.587 $Y2=2.815
r160 30 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.23 $Y=0.855
+ $X2=12.065 $Y2=0.855
r161 29 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.175 $Y=0.855
+ $X2=13.26 $Y2=0.94
r162 29 30 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=13.175 $Y=0.855
+ $X2=12.23 $Y2=0.855
r163 25 44 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.065 $Y=0.77
+ $X2=12.065 $Y2=0.855
r164 25 27 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=12.065 $Y=0.77
+ $X2=12.065 $Y2=0.515
r165 21 24 41.3382 $w=1.5e-07 $l=2.68e-07 $layer=POLY_cond $X=14.865 $Y=1.765
+ $X2=14.865 $Y2=1.497
r166 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.865 $Y=1.765
+ $X2=14.865 $Y2=2.4
r167 18 24 41.3382 $w=1.5e-07 $l=2.67e-07 $layer=POLY_cond $X=14.865 $Y=1.23
+ $X2=14.865 $Y2=1.497
r168 18 20 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=14.865 $Y=1.23
+ $X2=14.865 $Y2=0.74
r169 17 56 10.5996 $w=4.32e-07 $l=1.27279e-07 $layer=POLY_cond $X=13.985
+ $Y=1.425 $X2=13.895 $Y2=1.335
r170 16 24 6.9036 $w=3.9e-07 $l=1.20748e-07 $layer=POLY_cond $X=14.775 $Y=1.425
+ $X2=14.865 $Y2=1.497
r171 16 17 112.657 $w=3.9e-07 $l=7.9e-07 $layer=POLY_cond $X=14.775 $Y=1.425
+ $X2=13.985 $Y2=1.425
r172 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=13.895 $Y=2.245
+ $X2=13.895 $Y2=2.64
r173 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=13.895 $Y=2.155
+ $X2=13.895 $Y2=2.245
r174 11 56 23.3057 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=13.895 $Y=1.62
+ $X2=13.895 $Y2=1.335
r175 11 12 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=13.895 $Y=1.62
+ $X2=13.895 $Y2=2.155
r176 7 55 27.7542 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.875 $Y=1.05
+ $X2=13.875 $Y2=1.335
r177 7 9 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=13.875 $Y=1.05 $X2=13.875
+ $Y2=0.58
r178 2 47 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=12.305
+ $Y=1.96 $X2=12.455 $Y2=2.105
r179 2 33 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=12.305
+ $Y=1.96 $X2=12.455 $Y2=2.815
r180 1 44 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=11.925
+ $Y=0.37 $X2=12.065 $Y2=0.855
r181 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.925
+ $Y=0.37 $X2=12.065 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_27_74# 1 2 3 4 14 17 19 22 23 24 26 27
+ 28 31 35 38 42 44 47 49
r122 39 42 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.17 $Y=0.645
+ $X2=0.35 $Y2=0.645
r123 38 49 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.31 $Y=2.29
+ $X2=3.27 $Y2=2.375
r124 37 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=1.335
+ $X2=3.31 $Y2=1.25
r125 37 38 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.31 $Y=1.335
+ $X2=3.31 $Y2=2.29
r126 35 49 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=2.46 $X2=3.27
+ $Y2=2.375
r127 29 47 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.055 $Y=1.25
+ $X2=3.31 $Y2=1.25
r128 29 31 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.055 $Y=1.165
+ $X2=3.055 $Y2=0.765
r129 27 49 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.145 $Y=2.375
+ $X2=3.27 $Y2=2.375
r130 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.145 $Y=2.375
+ $X2=2.215 $Y2=2.375
r131 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=2.46
+ $X2=2.215 $Y2=2.375
r132 25 26 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.13 $Y=2.46
+ $X2=2.13 $Y2=2.905
r133 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=2.13 $Y2=2.905
r134 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=1.535 $Y2=2.99
r135 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.45 $Y=2.905
+ $X2=1.535 $Y2=2.99
r136 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.45 $Y=2.46
+ $X2=1.45 $Y2=2.905
r137 20 44 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.435 $Y=2.375
+ $X2=0.26 $Y2=2.375
r138 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.365 $Y=2.375
+ $X2=1.45 $Y2=2.46
r139 19 20 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.365 $Y=2.375
+ $X2=0.435 $Y2=2.375
r140 15 44 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.46
+ $X2=0.26 $Y2=2.375
r141 15 17 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=0.26 $Y=2.46
+ $X2=0.26 $Y2=2.465
r142 14 44 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.26 $Y2=2.375
r143 13 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=0.645
r144 13 14 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=2.29
r145 4 35 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.16
+ $Y=2.315 $X2=3.31 $Y2=2.46
r146 3 17 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.27 $Y2=2.465
r147 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.555 $X2=3.055 $Y2=0.765
r148 1 42 182 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.35 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 58 60 62 67 68 70 71 73 74 76 77 79 80 81 93 100 118 125 131 134 137 141
c161 3 0 9.53964e-20 $X=4.585 $Y=2.275
r162 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r163 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r164 134 135 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r165 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r166 129 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r167 129 138 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=13.68 $Y2=3.33
r168 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r169 126 137 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=13.785 $Y=3.33
+ $X2=13.557 $Y2=3.33
r170 126 128 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=13.785 $Y=3.33
+ $X2=14.64 $Y2=3.33
r171 125 140 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=15.005 $Y=3.33
+ $X2=15.182 $Y2=3.33
r172 125 128 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=15.005 $Y=3.33
+ $X2=14.64 $Y2=3.33
r173 124 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r174 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r175 121 124 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=13.2 $Y2=3.33
r176 120 123 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=13.2 $Y2=3.33
r177 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r178 118 137 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=13.33 $Y=3.33
+ $X2=13.557 $Y2=3.33
r179 118 123 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=13.33 $Y=3.33
+ $X2=13.2 $Y2=3.33
r180 117 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r181 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r182 114 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r183 113 114 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r184 111 114 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=9.84 $Y2=3.33
r185 110 113 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=9.84 $Y2=3.33
r186 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r187 108 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r188 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r189 105 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.49 $Y=3.33
+ $X2=6.325 $Y2=3.33
r190 105 107 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=6.49 $Y=3.33
+ $X2=7.44 $Y2=3.33
r191 104 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r192 104 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r193 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r194 101 131 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.13 $Y=3.33
+ $X2=5.005 $Y2=3.33
r195 101 103 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=5.13 $Y=3.33
+ $X2=6 $Y2=3.33
r196 100 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.16 $Y=3.33
+ $X2=6.325 $Y2=3.33
r197 100 103 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.16 $Y=3.33
+ $X2=6 $Y2=3.33
r198 99 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r199 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r200 96 99 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r201 95 98 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r202 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r203 93 131 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=5.005 $Y2=3.33
r204 93 98 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r205 92 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r206 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r207 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r208 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r209 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r210 85 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r212 81 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.92 $Y2=3.33
r213 81 108 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.44 $Y2=3.33
r214 79 116 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=10.8 $Y2=3.33
r215 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=11.07 $Y2=3.33
r216 78 120 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=11.235 $Y=3.33
+ $X2=11.28 $Y2=3.33
r217 78 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.235 $Y=3.33
+ $X2=11.07 $Y2=3.33
r218 76 113 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=9.865 $Y=3.33
+ $X2=9.84 $Y2=3.33
r219 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=3.33
+ $X2=10.03 $Y2=3.33
r220 75 116 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.8 $Y2=3.33
r221 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.03 $Y2=3.33
r222 73 107 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.51 $Y=3.33
+ $X2=7.44 $Y2=3.33
r223 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.51 $Y=3.33
+ $X2=7.675 $Y2=3.33
r224 72 110 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.84 $Y=3.33
+ $X2=7.92 $Y2=3.33
r225 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.84 $Y=3.33
+ $X2=7.675 $Y2=3.33
r226 70 91 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.16 $Y2=3.33
r227 70 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.51 $Y2=3.33
r228 69 95 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.64 $Y2=3.33
r229 69 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.51 $Y2=3.33
r230 67 84 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.72 $Y2=3.33
r231 67 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.07 $Y2=3.33
r232 66 88 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.2 $Y2=3.33
r233 66 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.07 $Y2=3.33
r234 62 65 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=15.13 $Y=1.985
+ $X2=15.13 $Y2=2.815
r235 60 140 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=15.13 $Y=3.245
+ $X2=15.182 $Y2=3.33
r236 60 65 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.13 $Y=3.245
+ $X2=15.13 $Y2=2.815
r237 56 137 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=13.557 $Y=3.245
+ $X2=13.557 $Y2=3.33
r238 56 58 11.3036 $w=4.53e-07 $l=4.3e-07 $layer=LI1_cond $X=13.557 $Y=3.245
+ $X2=13.557 $Y2=2.815
r239 52 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=3.245
+ $X2=11.07 $Y2=3.33
r240 52 54 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.07 $Y=3.245
+ $X2=11.07 $Y2=2.815
r241 48 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.03 $Y=3.245
+ $X2=10.03 $Y2=3.33
r242 48 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.03 $Y=3.245
+ $X2=10.03 $Y2=2.815
r243 44 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.675 $Y=3.245
+ $X2=7.675 $Y2=3.33
r244 44 46 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=7.675 $Y=3.245
+ $X2=7.675 $Y2=2.785
r245 40 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.325 $Y=3.245
+ $X2=6.325 $Y2=3.33
r246 40 42 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.325 $Y=3.245
+ $X2=6.325 $Y2=2.755
r247 36 131 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=3.33
r248 36 38 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=2.765
r249 32 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=3.33
r250 32 34 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=2.8
r251 28 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r252 28 30 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.805
r253 9 65 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.94
+ $Y=1.84 $X2=15.09 $Y2=2.815
r254 9 62 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.94
+ $Y=1.84 $X2=15.09 $Y2=1.985
r255 8 58 600 $w=1.7e-07 $l=4.10061e-07 $layer=licon1_PDIFF $count=1 $X=13.26
+ $Y=2.54 $X2=13.555 $Y2=2.815
r256 7 54 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=10.945
+ $Y=1.96 $X2=11.07 $Y2=2.815
r257 6 50 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.88
+ $Y=2.54 $X2=10.03 $Y2=2.815
r258 5 46 600 $w=1.7e-07 $l=1.00556e-06 $layer=licon1_PDIFF $count=1 $X=7.55
+ $Y=1.84 $X2=7.675 $Y2=2.785
r259 4 42 600 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=6.2
+ $Y=1.78 $X2=6.325 $Y2=2.755
r260 3 38 600 $w=1.7e-07 $l=6.52917e-07 $layer=licon1_PDIFF $count=1 $X=4.585
+ $Y=2.275 $X2=4.965 $Y2=2.765
r261 2 34 600 $w=1.7e-07 $l=6.47708e-07 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=2.315 $X2=2.47 $Y2=2.8
r262 1 30 600 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=1 $X=0.96
+ $Y=2.32 $X2=1.11 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%A_669_111# 1 2 3 4 5 6 21 24 25 26 28 30
+ 33 37 38 40 41 44 45 46 47 51 54 55 57 60 63 65 66 68 69
c194 63 0 1.85697e-19 $X=3.705 $Y=2.295
c195 57 0 7.11901e-20 $X=8.65 $Y=2.815
c196 37 0 1.64952e-19 $X=5.99 $Y=1.16
c197 25 0 9.53964e-20 $X=4.54 $Y=2.99
r198 65 66 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.805 $Y=2.377
+ $X2=5.64 $Y2=2.377
r199 62 63 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=3.65 $Y=0.995
+ $X2=3.65 $Y2=2.295
r200 60 62 10.6507 $w=3.43e-07 $l=2.3e-07 $layer=LI1_cond $X=3.562 $Y=0.765
+ $X2=3.562 $Y2=0.995
r201 55 57 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=8.18 $Y=2.855
+ $X2=8.65 $Y2=2.855
r202 54 55 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.095 $Y=2.73
+ $X2=8.18 $Y2=2.855
r203 53 54 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.095 $Y=2.5
+ $X2=8.095 $Y2=2.73
r204 49 51 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=8.11 $Y=1.48
+ $X2=8.11 $Y2=0.76
r205 48 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.79 $Y=2.415
+ $X2=7.705 $Y2=2.415
r206 47 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.01 $Y=2.415
+ $X2=8.095 $Y2=2.5
r207 47 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.01 $Y=2.415
+ $X2=7.79 $Y2=2.415
r208 45 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.985 $Y=1.565
+ $X2=8.11 $Y2=1.48
r209 45 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.985 $Y=1.565
+ $X2=7.79 $Y2=1.565
r210 44 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.705 $Y=2.33
+ $X2=7.705 $Y2=2.415
r211 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.705 $Y=1.65
+ $X2=7.79 $Y2=1.565
r212 43 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.705 $Y=1.65
+ $X2=7.705 $Y2=2.33
r213 41 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.62 $Y=2.415
+ $X2=7.705 $Y2=2.415
r214 41 68 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=7.62 $Y=2.415
+ $X2=6.16 $Y2=2.415
r215 40 68 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=2.377
+ $X2=6.16 $Y2=2.377
r216 40 65 12.7004 $w=2.43e-07 $l=2.7e-07 $layer=LI1_cond $X=6.075 $Y=2.377
+ $X2=5.805 $Y2=2.377
r217 39 40 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=6.075 $Y=1.245
+ $X2=6.075 $Y2=2.255
r218 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.99 $Y=1.16
+ $X2=6.075 $Y2=1.245
r219 37 38 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.99 $Y=1.16
+ $X2=5.795 $Y2=1.16
r220 31 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.63 $Y=1.075
+ $X2=5.795 $Y2=1.16
r221 31 33 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.63 $Y=1.075
+ $X2=5.63 $Y2=0.835
r222 30 66 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=4.71 $Y=2.34
+ $X2=5.64 $Y2=2.34
r223 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.625 $Y=2.425
+ $X2=4.71 $Y2=2.34
r224 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.625 $Y=2.425
+ $X2=4.625 $Y2=2.905
r225 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.54 $Y=2.99
+ $X2=4.625 $Y2=2.905
r226 25 26 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.54 $Y=2.99
+ $X2=3.845 $Y2=2.99
r227 22 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.705 $Y=2.905
+ $X2=3.845 $Y2=2.99
r228 22 24 18.3156 $w=2.78e-07 $l=4.45e-07 $layer=LI1_cond $X=3.705 $Y=2.905
+ $X2=3.705 $Y2=2.46
r229 21 63 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.705 $Y=2.435
+ $X2=3.705 $Y2=2.295
r230 21 24 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.705 $Y=2.435
+ $X2=3.705 $Y2=2.46
r231 6 57 600 $w=1.7e-07 $l=3.33729e-07 $layer=licon1_PDIFF $count=1 $X=8.52
+ $Y=2.54 $X2=8.65 $Y2=2.815
r232 5 65 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=5.655
+ $Y=2.275 $X2=5.805 $Y2=2.42
r233 4 24 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.61
+ $Y=2.315 $X2=3.76 $Y2=2.46
r234 3 51 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=8.01
+ $Y=0.485 $X2=8.15 $Y2=0.76
r235 2 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.49
+ $Y=0.625 $X2=5.63 $Y2=0.835
r236 1 60 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.345
+ $Y=0.555 $X2=3.555 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%Q 1 2 7 8 9 10 11 12 13
r19 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=14.645 $Y=2.405
+ $X2=14.645 $Y2=2.775
r20 11 12 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=14.645 $Y=1.985
+ $X2=14.645 $Y2=2.405
r21 10 11 10.8465 $w=3.38e-07 $l=3.2e-07 $layer=LI1_cond $X=14.645 $Y=1.665
+ $X2=14.645 $Y2=1.985
r22 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=14.645 $Y=1.295
+ $X2=14.645 $Y2=1.665
r23 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=14.645 $Y=0.925
+ $X2=14.645 $Y2=1.295
r24 7 8 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=14.645 $Y=0.515
+ $X2=14.645 $Y2=0.925
r25 2 13 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=14.515
+ $Y=1.84 $X2=14.64 $Y2=2.815
r26 2 11 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=14.515
+ $Y=1.84 $X2=14.64 $Y2=1.985
r27 1 7 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=14.505
+ $Y=0.37 $X2=14.65 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SEDFXTP_1%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 56 58 61 62 64 65 67 68 69 71 76 97 104 117 123 126 129 132 137 143 146
c173 30 0 1.72336e-19 $X=1.245 $Y=0.58
r174 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r175 141 143 9.13714 $w=6.83e-07 $l=7.5e-08 $layer=LI1_cond $X=13.68 $Y=0.257
+ $X2=13.755 $Y2=0.257
r176 141 142 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r177 139 141 1.57149 $w=6.83e-07 $l=9e-08 $layer=LI1_cond $X=13.59 $Y=0.257
+ $X2=13.68 $Y2=0.257
r178 136 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r179 135 139 6.80979 $w=6.83e-07 $l=3.9e-07 $layer=LI1_cond $X=13.2 $Y=0.257
+ $X2=13.59 $Y2=0.257
r180 135 137 14.812 $w=6.83e-07 $l=4e-07 $layer=LI1_cond $X=13.2 $Y=0.257
+ $X2=12.8 $Y2=0.257
r181 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r182 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r183 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r184 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r185 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r186 121 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r187 121 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=13.68 $Y2=0
r188 120 143 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=14.64 $Y=0
+ $X2=13.755 $Y2=0
r189 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r190 117 145 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=14.995 $Y=0
+ $X2=15.177 $Y2=0
r191 117 120 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.995 $Y=0
+ $X2=14.64 $Y2=0
r192 116 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r193 115 137 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=12.72 $Y=0 $X2=12.8
+ $Y2=0
r194 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r195 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r196 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r197 112 115 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r198 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r199 110 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.44 $Y=0
+ $X2=11.315 $Y2=0
r200 110 112 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.44 $Y=0
+ $X2=11.76 $Y2=0
r201 108 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r202 108 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=9.84 $Y2=0
r203 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r204 105 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10 $Y=0 $X2=9.875
+ $Y2=0
r205 105 107 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=10 $Y=0 $X2=10.8
+ $Y2=0
r206 104 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.19 $Y=0
+ $X2=11.315 $Y2=0
r207 104 107 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.19 $Y=0
+ $X2=10.8 $Y2=0
r208 103 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r209 102 103 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r210 99 102 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.44 $Y=0
+ $X2=9.36 $Y2=0
r211 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r212 97 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.75 $Y=0
+ $X2=9.875 $Y2=0
r213 97 102 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.75 $Y=0 $X2=9.36
+ $Y2=0
r214 96 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r215 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r216 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r217 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r218 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r219 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r220 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r221 87 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r222 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r223 84 87 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r224 84 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r225 83 86 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r226 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r227 81 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.235
+ $Y2=0
r228 81 83 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r229 80 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r230 80 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r231 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r232 77 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0
+ $X2=1.245 $Y2=0
r233 77 79 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.68
+ $Y2=0
r234 76 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0
+ $X2=2.235 $Y2=0
r235 76 79 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.68
+ $Y2=0
r236 74 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r237 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r238 71 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=0
+ $X2=1.245 $Y2=0
r239 71 73 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=0.72
+ $Y2=0
r240 69 103 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=9.36 $Y2=0
r241 69 100 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=7.44 $Y2=0
r242 67 95 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.005 $Y=0 $X2=6.96
+ $Y2=0
r243 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0 $X2=7.17
+ $Y2=0
r244 66 99 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=7.44 $Y2=0
r245 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.17
+ $Y2=0
r246 64 92 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.02 $Y=0 $X2=6 $Y2=0
r247 64 65 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.02 $Y=0 $X2=6.15
+ $Y2=0
r248 63 95 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.28 $Y=0 $X2=6.96
+ $Y2=0
r249 63 65 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.28 $Y=0 $X2=6.15
+ $Y2=0
r250 61 86 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=4.56 $Y2=0
r251 61 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.88
+ $Y2=0
r252 60 89 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.005 $Y=0 $X2=5.04
+ $Y2=0
r253 60 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.005 $Y=0 $X2=4.88
+ $Y2=0
r254 56 145 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=15.12 $Y=0.085
+ $X2=15.177 $Y2=0
r255 56 58 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.12 $Y=0.085
+ $X2=15.12 $Y2=0.515
r256 52 132 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.315 $Y=0.085
+ $X2=11.315 $Y2=0
r257 52 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.315 $Y=0.085
+ $X2=11.315 $Y2=0.515
r258 48 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.875 $Y=0.085
+ $X2=9.875 $Y2=0
r259 48 50 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.875 $Y=0.085
+ $X2=9.875 $Y2=0.515
r260 44 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.17 $Y=0.085
+ $X2=7.17 $Y2=0
r261 44 46 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.17 $Y=0.085
+ $X2=7.17 $Y2=0.55
r262 40 65 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0
r263 40 42 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0.665
r264 36 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0
r265 36 38 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0.805
r266 32 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0
r267 32 34 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0.765
r268 28 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r269 28 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.58
r270 9 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.94
+ $Y=0.37 $X2=15.08 $Y2=0.515
r271 8 139 91 $w=1.7e-07 $l=8.34356e-07 $layer=licon1_NDIFF $count=2 $X=12.825
+ $Y=0.37 $X2=13.59 $Y2=0.515
r272 7 54 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.13
+ $Y=0.37 $X2=11.275 $Y2=0.515
r273 6 50 182 $w=1.7e-07 $l=2.2951e-07 $layer=licon1_NDIFF $count=1 $X=9.7
+ $Y=0.485 $X2=9.915 $Y2=0.515
r274 5 46 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=7.025
+ $Y=0.37 $X2=7.17 $Y2=0.55
r275 4 42 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.37 $X2=6.185 $Y2=0.665
r276 3 38 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.7 $Y=0.625
+ $X2=4.84 $Y2=0.805
r277 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.095
+ $Y=0.555 $X2=2.235 $Y2=0.765
r278 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.37 $X2=1.245 $Y2=0.58
.ends

