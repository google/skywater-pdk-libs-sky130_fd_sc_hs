* File: sky130_fd_sc_hs__a2bb2o_1.pxi.spice
* Created: Thu Aug 27 20:27:38 2020
* 
x_PM_SKY130_FD_SC_HS__A2BB2O_1%A_93_264# N_A_93_264#_M1001_d N_A_93_264#_M1005_s
+ N_A_93_264#_c_81_n N_A_93_264#_M1002_g N_A_93_264#_M1008_g N_A_93_264#_c_83_n
+ N_A_93_264#_c_89_n N_A_93_264#_c_149_p N_A_93_264#_c_168_p N_A_93_264#_c_90_n
+ N_A_93_264#_c_91_n N_A_93_264#_c_92_n N_A_93_264#_c_84_n N_A_93_264#_c_94_n
+ N_A_93_264#_c_85_n N_A_93_264#_c_123_p N_A_93_264#_c_86_n N_A_93_264#_c_95_n
+ PM_SKY130_FD_SC_HS__A2BB2O_1%A_93_264#
x_PM_SKY130_FD_SC_HS__A2BB2O_1%A1_N N_A1_N_c_182_n N_A1_N_M1006_g N_A1_N_c_187_n
+ N_A1_N_M1003_g A1_N N_A1_N_c_184_n N_A1_N_c_185_n
+ PM_SKY130_FD_SC_HS__A2BB2O_1%A1_N
x_PM_SKY130_FD_SC_HS__A2BB2O_1%A2_N N_A2_N_c_224_n N_A2_N_M1011_g N_A2_N_c_225_n
+ N_A2_N_M1007_g A2_N PM_SKY130_FD_SC_HS__A2BB2O_1%A2_N
x_PM_SKY130_FD_SC_HS__A2BB2O_1%A_257_126# N_A_257_126#_M1006_d
+ N_A_257_126#_M1011_d N_A_257_126#_M1001_g N_A_257_126#_c_264_n
+ N_A_257_126#_M1005_g N_A_257_126#_c_265_n N_A_257_126#_c_266_n
+ N_A_257_126#_c_267_n N_A_257_126#_c_268_n N_A_257_126#_c_271_n
+ N_A_257_126#_c_272_n N_A_257_126#_c_273_n N_A_257_126#_c_269_n
+ PM_SKY130_FD_SC_HS__A2BB2O_1%A_257_126#
x_PM_SKY130_FD_SC_HS__A2BB2O_1%B2 N_B2_M1004_g N_B2_c_335_n N_B2_M1009_g B2
+ PM_SKY130_FD_SC_HS__A2BB2O_1%B2
x_PM_SKY130_FD_SC_HS__A2BB2O_1%B1 N_B1_M1010_g N_B1_c_371_n N_B1_c_372_n
+ N_B1_c_376_n N_B1_M1000_g B1 B1 N_B1_c_374_n PM_SKY130_FD_SC_HS__A2BB2O_1%B1
x_PM_SKY130_FD_SC_HS__A2BB2O_1%X N_X_M1008_s N_X_M1002_s N_X_c_401_n N_X_c_402_n
+ X X X N_X_c_405_n N_X_c_403_n X PM_SKY130_FD_SC_HS__A2BB2O_1%X
x_PM_SKY130_FD_SC_HS__A2BB2O_1%VPWR N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_c_424_n
+ N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n VPWR N_VPWR_c_428_n
+ N_VPWR_c_429_n N_VPWR_c_423_n N_VPWR_c_431_n PM_SKY130_FD_SC_HS__A2BB2O_1%VPWR
x_PM_SKY130_FD_SC_HS__A2BB2O_1%A_530_392# N_A_530_392#_M1005_d
+ N_A_530_392#_M1000_d N_A_530_392#_c_471_n N_A_530_392#_c_472_n
+ N_A_530_392#_c_473_n N_A_530_392#_c_474_n N_A_530_392#_c_475_n
+ PM_SKY130_FD_SC_HS__A2BB2O_1%A_530_392#
x_PM_SKY130_FD_SC_HS__A2BB2O_1%VGND N_VGND_M1008_d N_VGND_M1007_d N_VGND_M1010_d
+ N_VGND_c_501_n N_VGND_c_517_n N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_560_n
+ N_VGND_c_551_n N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n
+ N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n VGND N_VGND_c_511_n
+ N_VGND_c_512_n PM_SKY130_FD_SC_HS__A2BB2O_1%VGND
cc_1 VNB N_A_93_264#_c_81_n 0.0359931f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.765
cc_2 VNB N_A_93_264#_M1008_g 0.024394f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_3 VNB N_A_93_264#_c_83_n 3.96917e-19 $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.79
cc_4 VNB N_A_93_264#_c_84_n 0.00914112f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=1.79
cc_5 VNB N_A_93_264#_c_85_n 3.76316e-19 $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=1.12
cc_6 VNB N_A_93_264#_c_86_n 0.00668603f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.485
cc_7 VNB N_A1_N_c_182_n 0.00222805f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.96
cc_8 VNB A1_N 0.00271775f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.4
cc_9 VNB N_A1_N_c_184_n 0.0312696f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_10 VNB N_A1_N_c_185_n 0.0166691f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.65
cc_11 VNB N_A2_N_c_224_n 0.0384047f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=0.63
cc_12 VNB N_A2_N_c_225_n 0.0199265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A2_N 0.00300577f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.765
cc_14 VNB N_A_257_126#_M1001_g 0.020051f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.32
cc_15 VNB N_A_257_126#_c_264_n 0.0212895f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_16 VNB N_A_257_126#_c_265_n 0.00104163f $X=-0.19 $Y=-0.245 $X2=1.325
+ $Y2=1.875
cc_17 VNB N_A_257_126#_c_266_n 0.00564675f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.96
cc_18 VNB N_A_257_126#_c_267_n 0.0152508f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.875
cc_19 VNB N_A_257_126#_c_268_n 0.0462783f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.875
cc_20 VNB N_A_257_126#_c_269_n 0.00162172f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_21 VNB N_B2_M1004_g 0.0216081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B2_c_335_n 0.019829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB B2 0.00401095f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.4
cc_24 VNB N_B1_M1010_g 0.013239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_c_371_n 0.00886419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B1_c_372_n 0.0187569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB B1 0.0355701f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_28 VNB N_B1_c_374_n 0.0531247f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.96
cc_29 VNB N_X_c_401_n 0.02872f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.4
cc_30 VNB N_X_c_402_n 0.0124546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_403_n 0.0241894f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_32 VNB N_VPWR_c_423_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_33 VNB N_VGND_c_501_n 0.0122286f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_34 VNB N_VGND_c_502_n 0.00822066f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.905
cc_35 VNB N_VGND_c_503_n 0.0102407f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.875
cc_36 VNB N_VGND_c_504_n 0.0234937f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=1.79
cc_37 VNB N_VGND_c_505_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=2.905
cc_38 VNB N_VGND_c_506_n 0.0397362f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=2.635
cc_39 VNB N_VGND_c_507_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_508_n 0.00661898f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_41 VNB N_VGND_c_509_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_42 VNB N_VGND_c_510_n 0.022756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_511_n 0.0272571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_512_n 0.263154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A_93_264#_c_81_n 0.0273116f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.765
cc_46 VPB N_A_93_264#_c_83_n 0.00128976f $X=-0.19 $Y=1.66 $X2=0.815 $Y2=1.79
cc_47 VPB N_A_93_264#_c_89_n 0.00792166f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=1.875
cc_48 VPB N_A_93_264#_c_90_n 0.0156008f $X=-0.19 $Y=1.66 $X2=2.02 $Y2=1.875
cc_49 VPB N_A_93_264#_c_91_n 0.0119408f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=2.99
cc_50 VPB N_A_93_264#_c_92_n 0.00208946f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=2.99
cc_51 VPB N_A_93_264#_c_84_n 0.0028976f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=1.79
cc_52 VPB N_A_93_264#_c_94_n 0.0053202f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=2.635
cc_53 VPB N_A_93_264#_c_95_n 0.00661228f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.875
cc_54 VPB N_A1_N_c_182_n 0.00754378f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=1.96
cc_55 VPB N_A1_N_c_187_n 0.0203567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A2_N_c_224_n 0.0328712f $X=-0.19 $Y=1.66 $X2=2.595 $Y2=0.63
cc_57 VPB N_A_257_126#_c_264_n 0.0404586f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.81
cc_58 VPB N_A_257_126#_c_271_n 0.00773021f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=1.79
cc_59 VPB N_A_257_126#_c_272_n 0.00136291f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=2.635
cc_60 VPB N_A_257_126#_c_273_n 0.00592237f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=1.12
cc_61 VPB N_B2_c_335_n 0.0327973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB B2 0.00232698f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.4
cc_63 VPB N_B1_c_372_n 0.0112084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_B1_c_376_n 0.0287865f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.765
cc_65 VPB X 0.0481116f $X=-0.19 $Y=1.66 $X2=0.815 $Y2=1.65
cc_66 VPB N_X_c_405_n 0.0134975f $X=-0.19 $Y=1.66 $X2=2.735 $Y2=1.12
cc_67 VPB N_X_c_403_n 0.00770896f $X=-0.19 $Y=1.66 $X2=2.735 $Y2=1.12
cc_68 VPB N_VPWR_c_424_n 0.0062666f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.4
cc_69 VPB N_VPWR_c_425_n 0.00396743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_426_n 0.0227874f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=1.875
cc_71 VPB N_VPWR_c_427_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.9 $Y2=1.875
cc_72 VPB N_VPWR_c_428_n 0.0504791f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=1.21
cc_73 VPB N_VPWR_c_429_n 0.0278922f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=1.12
cc_74 VPB N_VPWR_c_423_n 0.0877203f $X=-0.19 $Y=1.66 $X2=2.735 $Y2=1.12
cc_75 VPB N_VPWR_c_431_n 0.00656574f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.485
cc_76 VPB N_A_530_392#_c_471_n 0.00663862f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.765
cc_77 VPB N_A_530_392#_c_472_n 0.00180901f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.4
cc_78 VPB N_A_530_392#_c_473_n 0.00856296f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.81
cc_79 VPB N_A_530_392#_c_474_n 0.0125972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_530_392#_c_475_n 0.0345863f $X=-0.19 $Y=1.66 $X2=0.815 $Y2=1.79
cc_81 N_A_93_264#_c_81_n N_A1_N_c_182_n 0.00867647f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_93_264#_c_83_n N_A1_N_c_182_n 0.00278959f $X=0.815 $Y=1.79 $X2=0 $Y2=0
cc_83 N_A_93_264#_c_89_n N_A1_N_c_182_n 0.0025073f $X=1.325 $Y=1.875 $X2=0 $Y2=0
cc_84 N_A_93_264#_c_86_n N_A1_N_c_182_n 6.91159e-19 $X=0.815 $Y=1.485 $X2=0
+ $Y2=0
cc_85 N_A_93_264#_c_81_n N_A1_N_c_187_n 0.0226094f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_93_264#_c_89_n N_A1_N_c_187_n 0.013516f $X=1.325 $Y=1.875 $X2=0 $Y2=0
cc_87 N_A_93_264#_c_92_n N_A1_N_c_187_n 0.00126785f $X=1.495 $Y=2.99 $X2=0 $Y2=0
cc_88 N_A_93_264#_c_81_n A1_N 2.74196e-19 $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_93_264#_M1008_g A1_N 0.00242144f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_90 N_A_93_264#_c_89_n A1_N 0.0189017f $X=1.325 $Y=1.875 $X2=0 $Y2=0
cc_91 N_A_93_264#_c_86_n A1_N 0.0239351f $X=0.815 $Y=1.485 $X2=0 $Y2=0
cc_92 N_A_93_264#_c_95_n A1_N 7.77974e-19 $X=1.41 $Y=1.875 $X2=0 $Y2=0
cc_93 N_A_93_264#_M1008_g N_A1_N_c_184_n 0.0205191f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_94 N_A_93_264#_c_89_n N_A1_N_c_184_n 0.00299885f $X=1.325 $Y=1.875 $X2=0
+ $Y2=0
cc_95 N_A_93_264#_c_86_n N_A1_N_c_184_n 0.00197815f $X=0.815 $Y=1.485 $X2=0
+ $Y2=0
cc_96 N_A_93_264#_M1008_g N_A1_N_c_185_n 0.0144354f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_97 N_A_93_264#_c_90_n N_A2_N_c_224_n 0.0198312f $X=2.02 $Y=1.875 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_93_264#_c_91_n N_A2_N_c_224_n 0.0146656f $X=2.185 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_93_264#_c_84_n N_A2_N_c_224_n 0.00653657f $X=2.105 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_93_264#_c_94_n N_A2_N_c_224_n 0.00311654f $X=2.35 $Y=2.635 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_93_264#_c_84_n N_A2_N_c_225_n 4.03823e-19 $X=2.105 $Y=1.79 $X2=0
+ $Y2=0
cc_102 N_A_93_264#_c_85_n N_A2_N_c_225_n 0.00551149f $X=2.19 $Y=1.12 $X2=0 $Y2=0
cc_103 N_A_93_264#_c_90_n A2_N 0.022839f $X=2.02 $Y=1.875 $X2=0 $Y2=0
cc_104 N_A_93_264#_c_84_n A2_N 0.0309176f $X=2.105 $Y=1.79 $X2=0 $Y2=0
cc_105 N_A_93_264#_c_85_n A2_N 0.00263878f $X=2.19 $Y=1.12 $X2=0 $Y2=0
cc_106 N_A_93_264#_c_91_n N_A_257_126#_M1011_d 0.00260133f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_107 N_A_93_264#_c_84_n N_A_257_126#_M1001_g 0.00584824f $X=2.105 $Y=1.79
+ $X2=0 $Y2=0
cc_108 N_A_93_264#_c_123_p N_A_257_126#_M1001_g 0.0108693f $X=2.735 $Y=1.12
+ $X2=0 $Y2=0
cc_109 N_A_93_264#_c_90_n N_A_257_126#_c_264_n 9.84486e-19 $X=2.02 $Y=1.875
+ $X2=0 $Y2=0
cc_110 N_A_93_264#_c_91_n N_A_257_126#_c_264_n 0.00661416f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_111 N_A_93_264#_c_84_n N_A_257_126#_c_264_n 0.00325837f $X=2.105 $Y=1.79
+ $X2=0 $Y2=0
cc_112 N_A_93_264#_c_94_n N_A_257_126#_c_264_n 0.00644697f $X=2.35 $Y=2.635
+ $X2=0 $Y2=0
cc_113 N_A_93_264#_c_123_p N_A_257_126#_c_264_n 0.00161323f $X=2.735 $Y=1.12
+ $X2=0 $Y2=0
cc_114 N_A_93_264#_M1008_g N_A_257_126#_c_266_n 6.54731e-19 $X=0.72 $Y=0.81
+ $X2=0 $Y2=0
cc_115 N_A_93_264#_M1005_s N_A_257_126#_c_271_n 0.0077352f $X=2.225 $Y=1.96
+ $X2=0 $Y2=0
cc_116 N_A_93_264#_c_90_n N_A_257_126#_c_271_n 0.0160722f $X=2.02 $Y=1.875 $X2=0
+ $Y2=0
cc_117 N_A_93_264#_c_91_n N_A_257_126#_c_271_n 0.00588659f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_118 N_A_93_264#_c_94_n N_A_257_126#_c_271_n 0.0226122f $X=2.35 $Y=2.635 $X2=0
+ $Y2=0
cc_119 N_A_93_264#_M1005_s N_A_257_126#_c_272_n 0.00301662f $X=2.225 $Y=1.96
+ $X2=0 $Y2=0
cc_120 N_A_93_264#_c_90_n N_A_257_126#_c_272_n 0.0143571f $X=2.02 $Y=1.875 $X2=0
+ $Y2=0
cc_121 N_A_93_264#_c_90_n N_A_257_126#_c_273_n 0.0244508f $X=2.02 $Y=1.875 $X2=0
+ $Y2=0
cc_122 N_A_93_264#_c_91_n N_A_257_126#_c_273_n 0.0204493f $X=2.185 $Y=2.99 $X2=0
+ $Y2=0
cc_123 N_A_93_264#_c_94_n N_A_257_126#_c_273_n 0.0204057f $X=2.35 $Y=2.635 $X2=0
+ $Y2=0
cc_124 N_A_93_264#_c_84_n N_A_257_126#_c_269_n 0.02533f $X=2.105 $Y=1.79 $X2=0
+ $Y2=0
cc_125 N_A_93_264#_c_123_p N_A_257_126#_c_269_n 0.0142216f $X=2.735 $Y=1.12
+ $X2=0 $Y2=0
cc_126 N_A_93_264#_c_123_p N_B2_M1004_g 0.00425018f $X=2.735 $Y=1.12 $X2=0 $Y2=0
cc_127 N_A_93_264#_c_91_n N_B2_c_335_n 3.01915e-19 $X=2.185 $Y=2.99 $X2=0 $Y2=0
cc_128 N_A_93_264#_c_123_p B2 0.00133508f $X=2.735 $Y=1.12 $X2=0 $Y2=0
cc_129 N_A_93_264#_c_123_p N_B1_M1010_g 5.52341e-19 $X=2.735 $Y=1.12 $X2=0 $Y2=0
cc_130 N_A_93_264#_M1008_g N_X_c_401_n 6.44746e-19 $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_131 N_A_93_264#_c_81_n N_X_c_402_n 0.00288561f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A_93_264#_c_86_n N_X_c_402_n 0.0101951f $X=0.815 $Y=1.485 $X2=0 $Y2=0
cc_133 N_A_93_264#_c_81_n N_X_c_405_n 0.0117704f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_93_264#_c_149_p N_X_c_405_n 0.0118053f $X=0.9 $Y=1.875 $X2=0 $Y2=0
cc_135 N_A_93_264#_c_86_n N_X_c_405_n 0.00792733f $X=0.815 $Y=1.485 $X2=0 $Y2=0
cc_136 N_A_93_264#_c_81_n N_X_c_403_n 0.0045674f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_93_264#_M1008_g N_X_c_403_n 0.00337861f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_138 N_A_93_264#_c_83_n N_X_c_403_n 0.0042417f $X=0.815 $Y=1.79 $X2=0 $Y2=0
cc_139 N_A_93_264#_c_86_n N_X_c_403_n 0.0253043f $X=0.815 $Y=1.485 $X2=0 $Y2=0
cc_140 N_A_93_264#_c_89_n N_VPWR_M1002_d 0.0015839f $X=1.325 $Y=1.875 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A_93_264#_c_149_p N_VPWR_M1002_d 7.23885e-19 $X=0.9 $Y=1.875 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_93_264#_c_81_n N_VPWR_c_424_n 0.0178031f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_93_264#_c_89_n N_VPWR_c_424_n 0.0151229f $X=1.325 $Y=1.875 $X2=0
+ $Y2=0
cc_144 N_A_93_264#_c_149_p N_VPWR_c_424_n 0.00687486f $X=0.9 $Y=1.875 $X2=0
+ $Y2=0
cc_145 N_A_93_264#_c_92_n N_VPWR_c_424_n 0.00802273f $X=1.495 $Y=2.99 $X2=0
+ $Y2=0
cc_146 N_A_93_264#_c_91_n N_VPWR_c_425_n 0.00280801f $X=2.185 $Y=2.99 $X2=0
+ $Y2=0
cc_147 N_A_93_264#_c_81_n N_VPWR_c_426_n 0.00413917f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_93_264#_c_91_n N_VPWR_c_428_n 0.0673515f $X=2.185 $Y=2.99 $X2=0 $Y2=0
cc_149 N_A_93_264#_c_92_n N_VPWR_c_428_n 0.0121867f $X=1.495 $Y=2.99 $X2=0 $Y2=0
cc_150 N_A_93_264#_c_81_n N_VPWR_c_423_n 0.00821711f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_93_264#_c_91_n N_VPWR_c_423_n 0.0379739f $X=2.185 $Y=2.99 $X2=0 $Y2=0
cc_152 N_A_93_264#_c_92_n N_VPWR_c_423_n 0.00660921f $X=1.495 $Y=2.99 $X2=0
+ $Y2=0
cc_153 N_A_93_264#_c_168_p A_258_392# 0.00412338f $X=1.41 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_93_264#_c_91_n N_A_530_392#_c_472_n 0.00522251f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_155 N_A_93_264#_c_94_n N_A_530_392#_c_472_n 0.0283016f $X=2.35 $Y=2.635 $X2=0
+ $Y2=0
cc_156 N_A_93_264#_c_85_n N_VGND_M1007_d 0.00555114f $X=2.19 $Y=1.12 $X2=0 $Y2=0
cc_157 N_A_93_264#_c_123_p N_VGND_M1007_d 0.00864797f $X=2.735 $Y=1.12 $X2=0
+ $Y2=0
cc_158 N_A_93_264#_M1008_g N_VGND_c_501_n 0.0147184f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_159 N_A_93_264#_c_86_n N_VGND_c_501_n 0.00542821f $X=0.815 $Y=1.485 $X2=0
+ $Y2=0
cc_160 N_A_93_264#_M1001_d N_VGND_c_517_n 0.00370806f $X=2.595 $Y=0.63 $X2=0
+ $Y2=0
cc_161 N_A_93_264#_c_85_n N_VGND_c_517_n 0.013831f $X=2.19 $Y=1.12 $X2=0 $Y2=0
cc_162 N_A_93_264#_c_123_p N_VGND_c_517_n 0.0389185f $X=2.735 $Y=1.12 $X2=0
+ $Y2=0
cc_163 N_A_93_264#_M1001_d N_VGND_c_502_n 6.84302e-19 $X=2.595 $Y=0.63 $X2=0
+ $Y2=0
cc_164 N_A_93_264#_M1008_g N_VGND_c_504_n 0.00438299f $X=0.72 $Y=0.81 $X2=0
+ $Y2=0
cc_165 N_A_93_264#_c_123_p N_VGND_c_510_n 0.00469776f $X=2.735 $Y=1.12 $X2=0
+ $Y2=0
cc_166 N_A_93_264#_M1008_g N_VGND_c_512_n 0.00439883f $X=0.72 $Y=0.81 $X2=0
+ $Y2=0
cc_167 N_A1_N_c_182_n N_A2_N_c_224_n 0.0162321f $X=1.215 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_168 N_A1_N_c_187_n N_A2_N_c_224_n 0.0541147f $X=1.215 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_169 A1_N N_A2_N_c_224_n 0.00115052f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_170 N_A1_N_c_184_n N_A2_N_c_224_n 0.0201104f $X=1.17 $Y=1.455 $X2=-0.19
+ $Y2=-0.245
cc_171 A1_N N_A2_N_c_225_n 3.7319e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_172 N_A1_N_c_185_n N_A2_N_c_225_n 0.0181059f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_173 A1_N A2_N 0.0281622f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A1_N_c_184_n A2_N 0.00114978f $X=1.17 $Y=1.455 $X2=0 $Y2=0
cc_175 N_A1_N_c_185_n A2_N 3.57707e-19 $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_176 A1_N N_A_257_126#_M1006_d 5.24173e-19 $X=1.115 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_177 N_A1_N_c_185_n N_A_257_126#_c_265_n 0.00103147f $X=1.17 $Y=1.29 $X2=0
+ $Y2=0
cc_178 N_A1_N_c_187_n N_VPWR_c_424_n 0.00594906f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_179 N_A1_N_c_187_n N_VPWR_c_428_n 0.00461464f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_180 N_A1_N_c_187_n N_VPWR_c_423_n 0.00908764f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_181 A1_N N_VGND_M1008_d 0.00184725f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_182 A1_N N_VGND_c_501_n 0.0014989f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A1_N_c_184_n N_VGND_c_501_n 0.0027243f $X=1.17 $Y=1.455 $X2=0 $Y2=0
cc_184 N_A1_N_c_185_n N_VGND_c_501_n 0.0031179f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_185 N_A1_N_c_185_n N_VGND_c_506_n 0.00412698f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_186 N_A1_N_c_185_n N_VGND_c_512_n 0.00468052f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_187 A2_N N_A_257_126#_M1006_d 2.07485e-19 $X=1.595 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A2_N_c_224_n N_A_257_126#_M1001_g 0.00209308f $X=1.605 $Y=1.885 $X2=0
+ $Y2=0
cc_189 N_A2_N_c_224_n N_A_257_126#_c_264_n 0.00502857f $X=1.605 $Y=1.885 $X2=0
+ $Y2=0
cc_190 N_A2_N_c_225_n N_A_257_126#_c_265_n 0.0172182f $X=1.64 $Y=1.29 $X2=0
+ $Y2=0
cc_191 A2_N N_A_257_126#_c_265_n 0.00272717f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A2_N_c_225_n N_A_257_126#_c_266_n 7.6083e-19 $X=1.64 $Y=1.29 $X2=0
+ $Y2=0
cc_193 N_A2_N_c_225_n N_A_257_126#_c_267_n 0.00657983f $X=1.64 $Y=1.29 $X2=0
+ $Y2=0
cc_194 A2_N N_A_257_126#_c_267_n 0.0044198f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_195 N_A2_N_c_225_n N_A_257_126#_c_268_n 3.36612e-19 $X=1.64 $Y=1.29 $X2=0
+ $Y2=0
cc_196 N_A2_N_c_224_n N_A_257_126#_c_272_n 0.00280662f $X=1.605 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_A2_N_c_224_n N_A_257_126#_c_273_n 0.00694327f $X=1.605 $Y=1.885 $X2=0
+ $Y2=0
cc_198 N_A2_N_c_224_n N_VPWR_c_428_n 0.00278271f $X=1.605 $Y=1.885 $X2=0 $Y2=0
cc_199 N_A2_N_c_224_n N_VPWR_c_423_n 0.00358137f $X=1.605 $Y=1.885 $X2=0 $Y2=0
cc_200 A2_N N_VGND_M1007_d 0.00228426f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_201 N_A2_N_c_224_n N_VGND_c_517_n 0.00115762f $X=1.605 $Y=1.885 $X2=0 $Y2=0
cc_202 A2_N N_VGND_c_517_n 0.0041082f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A2_N_c_225_n N_VGND_c_506_n 5.45085e-19 $X=1.64 $Y=1.29 $X2=0 $Y2=0
cc_204 N_A_257_126#_c_268_n N_B2_M1004_g 0.0270626f $X=2.43 $Y=0.355 $X2=0 $Y2=0
cc_205 N_A_257_126#_c_264_n N_B2_c_335_n 0.0338295f $X=2.575 $Y=1.885 $X2=0
+ $Y2=0
cc_206 N_A_257_126#_c_272_n N_B2_c_335_n 8.87777e-19 $X=2.445 $Y=2.13 $X2=0
+ $Y2=0
cc_207 N_A_257_126#_c_269_n N_B2_c_335_n 4.14706e-19 $X=2.5 $Y=1.615 $X2=0 $Y2=0
cc_208 N_A_257_126#_c_264_n B2 0.00114361f $X=2.575 $Y=1.885 $X2=0 $Y2=0
cc_209 N_A_257_126#_c_269_n B2 0.0208896f $X=2.5 $Y=1.615 $X2=0 $Y2=0
cc_210 N_A_257_126#_c_264_n N_VPWR_c_425_n 5.74104e-19 $X=2.575 $Y=1.885 $X2=0
+ $Y2=0
cc_211 N_A_257_126#_c_264_n N_VPWR_c_428_n 0.0044313f $X=2.575 $Y=1.885 $X2=0
+ $Y2=0
cc_212 N_A_257_126#_c_264_n N_VPWR_c_423_n 0.00859008f $X=2.575 $Y=1.885 $X2=0
+ $Y2=0
cc_213 N_A_257_126#_c_264_n N_A_530_392#_c_471_n 7.38235e-19 $X=2.575 $Y=1.885
+ $X2=0 $Y2=0
cc_214 N_A_257_126#_c_272_n N_A_530_392#_c_471_n 0.012587f $X=2.445 $Y=2.13
+ $X2=0 $Y2=0
cc_215 N_A_257_126#_c_264_n N_A_530_392#_c_472_n 0.00552396f $X=2.575 $Y=1.885
+ $X2=0 $Y2=0
cc_216 N_A_257_126#_c_271_n N_A_530_392#_c_472_n 0.0125099f $X=2.36 $Y=2.215
+ $X2=0 $Y2=0
cc_217 N_A_257_126#_c_272_n N_A_530_392#_c_472_n 5.91945e-19 $X=2.445 $Y=2.13
+ $X2=0 $Y2=0
cc_218 N_A_257_126#_c_265_n N_VGND_c_501_n 0.0223974f $X=1.425 $Y=0.845 $X2=0
+ $Y2=0
cc_219 N_A_257_126#_c_266_n N_VGND_c_501_n 0.0219867f $X=1.59 $Y=0.387 $X2=0
+ $Y2=0
cc_220 N_A_257_126#_M1001_g N_VGND_c_517_n 0.00837945f $X=2.52 $Y=0.95 $X2=0
+ $Y2=0
cc_221 N_A_257_126#_c_267_n N_VGND_c_517_n 0.0573731f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_222 N_A_257_126#_c_268_n N_VGND_c_517_n 0.00391065f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_223 N_A_257_126#_c_267_n N_VGND_c_502_n 0.0210179f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_224 N_A_257_126#_c_268_n N_VGND_c_502_n 0.00727503f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_225 N_A_257_126#_c_266_n N_VGND_c_506_n 0.0218645f $X=1.59 $Y=0.387 $X2=0
+ $Y2=0
cc_226 N_A_257_126#_c_267_n N_VGND_c_506_n 0.0657312f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_227 N_A_257_126#_c_268_n N_VGND_c_506_n 0.00641604f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_228 N_A_257_126#_c_266_n N_VGND_c_512_n 0.0118577f $X=1.59 $Y=0.387 $X2=0
+ $Y2=0
cc_229 N_A_257_126#_c_267_n N_VGND_c_512_n 0.0366452f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_230 N_A_257_126#_c_268_n N_VGND_c_512_n 0.00987452f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_231 N_B2_c_335_n N_B1_c_372_n 0.0249358f $X=3.025 $Y=1.885 $X2=0 $Y2=0
cc_232 B2 N_B1_c_372_n 0.00756601f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B2_c_335_n N_B1_c_376_n 0.0185501f $X=3.025 $Y=1.885 $X2=0 $Y2=0
cc_234 N_B2_M1004_g N_B1_c_374_n 0.0258771f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_235 N_B2_c_335_n N_VPWR_c_425_n 0.0111542f $X=3.025 $Y=1.885 $X2=0 $Y2=0
cc_236 N_B2_c_335_n N_VPWR_c_428_n 0.00413917f $X=3.025 $Y=1.885 $X2=0 $Y2=0
cc_237 N_B2_c_335_n N_VPWR_c_423_n 0.0081781f $X=3.025 $Y=1.885 $X2=0 $Y2=0
cc_238 N_B2_c_335_n N_A_530_392#_c_471_n 2.72398e-19 $X=3.025 $Y=1.885 $X2=0
+ $Y2=0
cc_239 B2 N_A_530_392#_c_471_n 8.43333e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_240 N_B2_c_335_n N_A_530_392#_c_472_n 0.00554978f $X=3.025 $Y=1.885 $X2=0
+ $Y2=0
cc_241 N_B2_c_335_n N_A_530_392#_c_473_n 0.0170729f $X=3.025 $Y=1.885 $X2=0
+ $Y2=0
cc_242 B2 N_A_530_392#_c_473_n 0.0258292f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_243 N_B2_M1004_g N_VGND_c_517_n 0.00564957f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_244 B2 N_VGND_c_517_n 9.81631e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_245 N_B2_M1004_g N_VGND_c_502_n 0.00515291f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_246 N_B2_M1004_g N_VGND_c_503_n 0.00266787f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_247 N_B2_M1004_g N_VGND_c_551_n 0.00425334f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_248 N_B2_c_335_n N_VGND_c_551_n 0.00117163f $X=3.025 $Y=1.885 $X2=0 $Y2=0
cc_249 B2 N_VGND_c_551_n 0.00366871f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_250 N_B2_M1004_g N_VGND_c_508_n 0.00246733f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_251 N_B2_M1004_g N_VGND_c_510_n 0.00102955f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_252 N_B2_M1004_g N_VGND_c_512_n 0.00283952f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_253 N_B1_c_376_n N_VPWR_c_425_n 0.0142316f $X=3.505 $Y=1.885 $X2=0 $Y2=0
cc_254 N_B1_c_376_n N_VPWR_c_429_n 0.00413917f $X=3.505 $Y=1.885 $X2=0 $Y2=0
cc_255 N_B1_c_376_n N_VPWR_c_423_n 0.00822528f $X=3.505 $Y=1.885 $X2=0 $Y2=0
cc_256 N_B1_c_376_n N_A_530_392#_c_473_n 0.0181223f $X=3.505 $Y=1.885 $X2=0
+ $Y2=0
cc_257 N_B1_c_376_n N_A_530_392#_c_474_n 4.02768e-19 $X=3.505 $Y=1.885 $X2=0
+ $Y2=0
cc_258 N_B1_c_376_n N_A_530_392#_c_475_n 0.00634858f $X=3.505 $Y=1.885 $X2=0
+ $Y2=0
cc_259 B1 N_VGND_M1010_d 0.0022726f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_260 B1 N_VGND_c_503_n 0.0330236f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_261 N_B1_c_374_n N_VGND_c_503_n 0.0137935f $X=3.65 $Y=0.355 $X2=0 $Y2=0
cc_262 N_B1_M1010_g N_VGND_c_560_n 0.0124674f $X=3.49 $Y=0.95 $X2=0 $Y2=0
cc_263 B1 N_VGND_c_560_n 0.00390864f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_264 N_B1_M1010_g N_VGND_c_510_n 0.00872234f $X=3.49 $Y=0.95 $X2=0 $Y2=0
cc_265 N_B1_c_371_n N_VGND_c_510_n 0.00112456f $X=3.505 $Y=1.435 $X2=0 $Y2=0
cc_266 B1 N_VGND_c_510_n 0.0221741f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_267 N_B1_c_374_n N_VGND_c_510_n 0.00120812f $X=3.65 $Y=0.355 $X2=0 $Y2=0
cc_268 B1 N_VGND_c_511_n 0.0476503f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_269 N_B1_c_374_n N_VGND_c_511_n 0.00865075f $X=3.65 $Y=0.355 $X2=0 $Y2=0
cc_270 B1 N_VGND_c_512_n 0.0257336f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_271 N_B1_c_374_n N_VGND_c_512_n 0.0119279f $X=3.65 $Y=0.355 $X2=0 $Y2=0
cc_272 X N_VPWR_c_424_n 0.0595244f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_273 X N_VPWR_c_426_n 0.0193209f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_274 X N_VPWR_c_423_n 0.0159921f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_275 N_X_c_401_n N_VGND_c_501_n 0.021946f $X=0.505 $Y=0.585 $X2=0 $Y2=0
cc_276 N_X_c_401_n N_VGND_c_504_n 0.0161045f $X=0.505 $Y=0.585 $X2=0 $Y2=0
cc_277 N_X_c_401_n N_VGND_c_512_n 0.0163598f $X=0.505 $Y=0.585 $X2=0 $Y2=0
cc_278 N_VPWR_c_425_n N_A_530_392#_c_472_n 0.0452765f $X=3.265 $Y=2.455 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_428_n N_A_530_392#_c_472_n 0.00749631f $X=3.085 $Y=3.33 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_423_n N_A_530_392#_c_472_n 0.0062048f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_281 N_VPWR_M1009_d N_A_530_392#_c_473_n 0.00229612f $X=3.1 $Y=1.96 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_425_n N_A_530_392#_c_473_n 0.0196221f $X=3.265 $Y=2.455 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_425_n N_A_530_392#_c_475_n 0.0465996f $X=3.265 $Y=2.455 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_429_n N_A_530_392#_c_475_n 0.011066f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_285 N_VPWR_c_423_n N_A_530_392#_c_475_n 0.00915947f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_286 N_A_530_392#_c_473_n N_VGND_c_510_n 0.00300932f $X=3.645 $Y=2.035 $X2=0
+ $Y2=0
cc_287 N_A_530_392#_c_474_n N_VGND_c_510_n 0.00793931f $X=3.77 $Y=2.12 $X2=0
+ $Y2=0
cc_288 N_VGND_c_503_n A_605_126# 0.00487694f $X=3.23 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_289 N_VGND_c_560_n A_605_126# 0.00244694f $X=3.54 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_290 N_VGND_c_551_n A_605_126# 0.00779459f $X=3.315 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
