# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.785000 2.025000 2.115000 2.355000 ;
        RECT 1.945000 1.125000 2.305000 1.780000 ;
        RECT 1.945000 1.780000 2.115000 2.025000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.116000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.800000 9.035000 1.970000 ;
        RECT 7.805000 1.970000 8.135000 2.980000 ;
        RECT 7.820000 0.350000 8.150000 0.960000 ;
        RECT 7.820000 0.960000 9.035000 1.130000 ;
        RECT 8.700000 0.350000 9.035000 0.960000 ;
        RECT 8.705000 1.970000 9.035000 2.980000 ;
        RECT 8.865000 1.130000 9.035000 1.800000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.505000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.960000 ;
      RECT 0.115000  0.960000 1.135000 1.130000 ;
      RECT 0.115000  1.950000 0.845000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.625000  0.085000 0.795000 0.790000 ;
      RECT 0.645000  2.290000 0.815000 3.245000 ;
      RECT 0.675000  1.130000 1.135000 1.550000 ;
      RECT 0.675000  1.550000 0.845000 1.950000 ;
      RECT 0.965000  0.255000 1.815000 0.425000 ;
      RECT 0.965000  0.425000 1.135000 0.960000 ;
      RECT 1.015000  1.820000 1.475000 2.525000 ;
      RECT 1.015000  2.525000 2.165000 2.695000 ;
      RECT 1.015000  2.695000 1.475000 2.980000 ;
      RECT 1.305000  0.595000 1.475000 1.220000 ;
      RECT 1.305000  1.220000 1.765000 1.550000 ;
      RECT 1.305000  1.550000 1.475000 1.820000 ;
      RECT 1.645000  0.425000 1.815000 0.730000 ;
      RECT 1.645000  0.730000 2.655000 0.900000 ;
      RECT 1.655000  2.865000 1.825000 3.245000 ;
      RECT 1.985000  0.085000 2.315000 0.560000 ;
      RECT 1.995000  2.695000 2.165000 2.905000 ;
      RECT 1.995000  2.905000 3.375000 3.075000 ;
      RECT 2.335000  1.950000 2.645000 2.120000 ;
      RECT 2.335000  2.120000 2.505000 2.735000 ;
      RECT 2.475000  1.070000 2.995000 1.240000 ;
      RECT 2.475000  1.240000 2.645000 1.950000 ;
      RECT 2.485000  0.255000 3.875000 0.425000 ;
      RECT 2.485000  0.425000 2.655000 0.730000 ;
      RECT 2.705000  2.485000 3.035000 2.735000 ;
      RECT 2.815000  1.410000 3.345000 1.580000 ;
      RECT 2.815000  1.580000 2.985000 2.250000 ;
      RECT 2.815000  2.250000 4.385000 2.420000 ;
      RECT 2.815000  2.420000 3.035000 2.485000 ;
      RECT 2.825000  0.595000 2.995000 1.070000 ;
      RECT 3.155000  1.750000 3.875000 2.080000 ;
      RECT 3.175000  0.620000 3.535000 0.950000 ;
      RECT 3.175000  0.950000 3.345000 1.410000 ;
      RECT 3.205000  2.590000 4.385000 2.760000 ;
      RECT 3.205000  2.760000 3.375000 2.905000 ;
      RECT 3.705000  0.425000 3.875000 0.690000 ;
      RECT 3.705000  0.690000 4.680000 0.860000 ;
      RECT 3.705000  0.860000 3.875000 1.750000 ;
      RECT 3.715000  2.930000 4.045000 3.245000 ;
      RECT 4.045000  1.030000 5.020000 1.200000 ;
      RECT 4.045000  1.200000 4.725000 1.370000 ;
      RECT 4.055000  1.630000 4.385000 2.250000 ;
      RECT 4.090000  0.085000 4.340000 0.520000 ;
      RECT 4.215000  2.760000 4.385000 2.905000 ;
      RECT 4.215000  2.905000 5.955000 3.075000 ;
      RECT 4.510000  0.255000 5.995000 0.425000 ;
      RECT 4.510000  0.425000 4.680000 0.690000 ;
      RECT 4.555000  1.370000 4.725000 2.735000 ;
      RECT 4.850000  0.595000 5.180000 0.950000 ;
      RECT 4.850000  0.950000 5.020000 1.030000 ;
      RECT 4.895000  1.370000 5.520000 1.540000 ;
      RECT 4.895000  1.540000 5.065000 2.905000 ;
      RECT 5.190000  1.150000 5.520000 1.370000 ;
      RECT 5.235000  1.710000 5.860000 1.880000 ;
      RECT 5.235000  1.880000 5.405000 2.735000 ;
      RECT 5.350000  0.720000 5.860000 0.970000 ;
      RECT 5.625000  2.050000 5.955000 2.905000 ;
      RECT 5.665000  0.425000 5.995000 0.510000 ;
      RECT 5.690000  0.970000 5.860000 1.140000 ;
      RECT 5.690000  1.140000 6.800000 1.220000 ;
      RECT 5.690000  1.220000 7.130000 1.310000 ;
      RECT 5.690000  1.310000 5.860000 1.710000 ;
      RECT 6.130000  1.480000 6.460000 1.720000 ;
      RECT 6.130000  1.720000 7.470000 1.810000 ;
      RECT 6.290000  1.810000 7.470000 1.890000 ;
      RECT 6.315000  2.450000 6.650000 3.245000 ;
      RECT 6.410000  0.085000 6.660000 0.970000 ;
      RECT 6.630000  1.310000 7.130000 1.390000 ;
      RECT 6.800000  1.390000 7.130000 1.550000 ;
      RECT 6.820000  1.890000 7.150000 2.980000 ;
      RECT 6.890000  0.350000 7.140000 0.880000 ;
      RECT 6.890000  0.880000 7.470000 0.970000 ;
      RECT 6.970000  0.970000 7.470000 1.050000 ;
      RECT 7.300000  1.050000 7.470000 1.300000 ;
      RECT 7.300000  1.300000 8.665000 1.630000 ;
      RECT 7.300000  1.630000 7.470000 1.720000 ;
      RECT 7.320000  0.085000 7.650000 0.710000 ;
      RECT 7.355000  2.060000 7.605000 3.245000 ;
      RECT 8.330000  0.085000 8.500000 0.790000 ;
      RECT 8.335000  2.140000 8.505000 3.245000 ;
      RECT 9.210000  0.085000 9.460000 1.130000 ;
      RECT 9.235000  1.820000 9.485000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_hs__dfxtp_4
