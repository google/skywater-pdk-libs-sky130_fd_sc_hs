* File: sky130_fd_sc_hs__a2111o_4.pex.spice
* Created: Tue Sep  1 19:48:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2111O_4%A_137_260# 1 2 3 4 5 16 18 19 21 24 26 28
+ 31 33 35 38 42 44 51 54 57 59 62 66 68 72 74 78 80 81 85 87 90
c182 87 0 7.64327e-20 $X=4.135 $Y=1.005
c183 81 0 1.34483e-19 $X=3.13 $Y=1.465
c184 78 0 1.83628e-19 $X=6.605 $Y=0.79
c185 74 0 7.29804e-20 $X=6.51 $Y=1.195
c186 72 0 8.41147e-20 $X=5.005 $Y=0.515
c187 66 0 1.39795e-19 $X=4.135 $Y=0.515
c188 59 0 1.80394e-19 $X=3.13 $Y=1.95
c189 54 0 1.47805e-19 $X=3.265 $Y=0.515
r190 97 98 2.54354 $w=3.79e-07 $l=2e-08 $layer=POLY_cond $X=2.125 $Y=1.532
+ $X2=2.145 $Y2=1.532
r191 96 97 52.1425 $w=3.79e-07 $l=4.1e-07 $layer=POLY_cond $X=1.715 $Y=1.532
+ $X2=2.125 $Y2=1.532
r192 95 96 5.08707 $w=3.79e-07 $l=4e-08 $layer=POLY_cond $X=1.675 $Y=1.532
+ $X2=1.715 $Y2=1.532
r193 94 95 49.5989 $w=3.79e-07 $l=3.9e-07 $layer=POLY_cond $X=1.285 $Y=1.532
+ $X2=1.675 $Y2=1.532
r194 93 94 7.63061 $w=3.79e-07 $l=6e-08 $layer=POLY_cond $X=1.225 $Y=1.532
+ $X2=1.285 $Y2=1.532
r195 87 88 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.135 $Y=1.005
+ $X2=4.135 $Y2=1.195
r196 82 85 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.13 $Y=2.035
+ $X2=3.32 $Y2=2.035
r197 76 78 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=6.64 $Y=1.11
+ $X2=6.64 $Y2=0.79
r198 75 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=1.195
+ $X2=5.005 $Y2=1.195
r199 74 76 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.51 $Y=1.195
+ $X2=6.64 $Y2=1.11
r200 74 75 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=6.51 $Y=1.195
+ $X2=5.09 $Y2=1.195
r201 70 90 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=1.11
+ $X2=5.005 $Y2=1.195
r202 70 72 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.005 $Y=1.11
+ $X2=5.005 $Y2=0.515
r203 69 88 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.22 $Y=1.195
+ $X2=4.135 $Y2=1.195
r204 68 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=1.195
+ $X2=5.005 $Y2=1.195
r205 68 69 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.92 $Y=1.195
+ $X2=4.22 $Y2=1.195
r206 64 87 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=0.92
+ $X2=4.135 $Y2=1.005
r207 64 66 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.135 $Y=0.92
+ $X2=4.135 $Y2=0.515
r208 63 80 2.57001 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.35 $Y=1.005
+ $X2=3.197 $Y2=1.005
r209 62 87 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=1.005
+ $X2=4.135 $Y2=1.005
r210 62 63 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.05 $Y=1.005
+ $X2=3.35 $Y2=1.005
r211 59 82 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=1.95
+ $X2=3.13 $Y2=2.035
r212 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=1.63
+ $X2=3.13 $Y2=1.465
r213 58 59 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.13 $Y=1.63
+ $X2=3.13 $Y2=1.95
r214 57 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=1.3
+ $X2=3.13 $Y2=1.465
r215 56 80 3.87901 $w=2.37e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.13 $Y=1.09
+ $X2=3.197 $Y2=1.005
r216 56 57 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.13 $Y=1.09
+ $X2=3.13 $Y2=1.3
r217 52 80 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=3.197 $Y=0.92
+ $X2=3.197 $Y2=1.005
r218 52 54 15.3029 $w=3.03e-07 $l=4.05e-07 $layer=LI1_cond $X=3.197 $Y=0.92
+ $X2=3.197 $Y2=0.515
r219 51 100 11.4459 $w=3.79e-07 $l=9e-08 $layer=POLY_cond $X=2.485 $Y=1.532
+ $X2=2.575 $Y2=1.532
r220 51 98 43.2401 $w=3.79e-07 $l=3.4e-07 $layer=POLY_cond $X=2.485 $Y=1.532
+ $X2=2.145 $Y2=1.532
r221 50 51 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.485
+ $Y=1.465 $X2=2.485 $Y2=1.465
r222 47 93 24.1636 $w=3.79e-07 $l=1.9e-07 $layer=POLY_cond $X=1.035 $Y=1.532
+ $X2=1.225 $Y2=1.532
r223 47 91 33.066 $w=3.79e-07 $l=2.6e-07 $layer=POLY_cond $X=1.035 $Y=1.532
+ $X2=0.775 $Y2=1.532
r224 46 50 50.6376 $w=3.28e-07 $l=1.45e-06 $layer=LI1_cond $X=1.035 $Y=1.465
+ $X2=2.485 $Y2=1.465
r225 46 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.035
+ $Y=1.465 $X2=1.035 $Y2=1.465
r226 44 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=1.465
+ $X2=3.13 $Y2=1.465
r227 44 50 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.045 $Y=1.465
+ $X2=2.485 $Y2=1.465
r228 40 100 24.5487 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.575 $Y=1.3
+ $X2=2.575 $Y2=1.532
r229 40 42 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.575 $Y=1.3
+ $X2=2.575 $Y2=0.74
r230 36 98 24.5487 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.145 $Y=1.3
+ $X2=2.145 $Y2=1.532
r231 36 38 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.145 $Y=1.3
+ $X2=2.145 $Y2=0.74
r232 33 97 24.5487 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.125 $Y=1.765
+ $X2=2.125 $Y2=1.532
r233 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.125 $Y=1.765
+ $X2=2.125 $Y2=2.4
r234 29 96 24.5487 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.715 $Y=1.3
+ $X2=1.715 $Y2=1.532
r235 29 31 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.715 $Y=1.3
+ $X2=1.715 $Y2=0.74
r236 26 95 24.5487 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.675 $Y=1.765
+ $X2=1.675 $Y2=1.532
r237 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.675 $Y=1.765
+ $X2=1.675 $Y2=2.4
r238 22 94 24.5487 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.285 $Y=1.3
+ $X2=1.285 $Y2=1.532
r239 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.285 $Y=1.3
+ $X2=1.285 $Y2=0.74
r240 19 93 24.5487 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.225 $Y=1.765
+ $X2=1.225 $Y2=1.532
r241 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.225 $Y=1.765
+ $X2=1.225 $Y2=2.4
r242 16 91 24.5487 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.775 $Y=1.765
+ $X2=0.775 $Y2=1.532
r243 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.775 $Y=1.765
+ $X2=0.775 $Y2=2.4
r244 5 85 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=3.17
+ $Y=1.96 $X2=3.32 $Y2=2.115
r245 4 78 182 $w=1.7e-07 $l=4.84974e-07 $layer=licon1_NDIFF $count=1 $X=6.465
+ $Y=0.37 $X2=6.605 $Y2=0.79
r246 3 72 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.865
+ $Y=0.37 $X2=5.005 $Y2=0.515
r247 2 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.995
+ $Y=0.37 $X2=4.135 $Y2=0.515
r248 1 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.125
+ $Y=0.37 $X2=3.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%D1 3 6 7 9 12 15 16 18 19 25 26
c67 15 0 1.34483e-19 $X=3.545 $Y=1.795
c68 12 0 1.47805e-19 $X=3.48 $Y=0.69
r69 26 27 9.76012 $w=3.21e-07 $l=6.5e-08 $layer=POLY_cond $X=3.48 $Y=1.425
+ $X2=3.545 $Y2=1.425
r70 24 26 1.50156 $w=3.21e-07 $l=1e-08 $layer=POLY_cond $X=3.47 $Y=1.425
+ $X2=3.48 $Y2=1.425
r71 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.425 $X2=3.47 $Y2=1.425
r72 22 24 56.3084 $w=3.21e-07 $l=3.75e-07 $layer=POLY_cond $X=3.095 $Y=1.425
+ $X2=3.47 $Y2=1.425
r73 21 22 6.75701 $w=3.21e-07 $l=4.5e-08 $layer=POLY_cond $X=3.05 $Y=1.425
+ $X2=3.095 $Y2=1.425
r74 19 25 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=1.425
r75 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.545 $Y=1.885
+ $X2=3.545 $Y2=2.46
r76 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.545 $Y=1.795
+ $X2=3.545 $Y2=1.885
r77 14 27 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.545 $Y=1.59
+ $X2=3.545 $Y2=1.425
r78 14 15 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.545 $Y=1.59
+ $X2=3.545 $Y2=1.795
r79 10 26 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.26
+ $X2=3.48 $Y2=1.425
r80 10 12 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.48 $Y=1.26
+ $X2=3.48 $Y2=0.69
r81 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.095 $Y=1.885
+ $X2=3.095 $Y2=2.46
r82 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.095 $Y=1.795 $X2=3.095
+ $Y2=1.885
r83 5 22 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=1.59
+ $X2=3.095 $Y2=1.425
r84 5 6 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.095 $Y=1.59
+ $X2=3.095 $Y2=1.795
r85 1 21 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.26
+ $X2=3.05 $Y2=1.425
r86 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.05 $Y=1.26 $X2=3.05
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%C1 3 5 7 10 12 13 15 16 17 18 19 20 27
c66 17 0 8.41147e-20 $X=4.36 $Y=1.235
c67 12 0 7.64327e-20 $X=4.37 $Y=1.45
c68 3 0 1.39795e-19 $X=3.92 $Y=0.69
r69 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.46
+ $Y=1.615 $X2=4.46 $Y2=1.615
r70 27 29 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=4.445 $Y=1.667
+ $X2=4.46 $Y2=1.667
r71 26 27 9.93132 $w=3.64e-07 $l=7.5e-08 $layer=POLY_cond $X=4.37 $Y=1.667
+ $X2=4.445 $Y2=1.667
r72 25 26 49.6566 $w=3.64e-07 $l=3.75e-07 $layer=POLY_cond $X=3.995 $Y=1.667
+ $X2=4.37 $Y2=1.667
r73 24 25 9.93132 $w=3.64e-07 $l=7.5e-08 $layer=POLY_cond $X=3.92 $Y=1.667
+ $X2=3.995 $Y2=1.667
r74 19 20 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=5.04 $Y2=1.615
r75 19 30 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=4.56 $Y=1.615 $X2=4.46
+ $Y2=1.615
r76 18 30 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=4.08 $Y=1.615
+ $X2=4.46 $Y2=1.615
r77 16 17 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=4.36 $Y=1.085
+ $X2=4.36 $Y2=1.235
r78 13 27 23.572 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=4.445 $Y=1.885
+ $X2=4.445 $Y2=1.667
r79 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.445 $Y=1.885
+ $X2=4.445 $Y2=2.46
r80 12 26 23.572 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=4.37 $Y=1.45
+ $X2=4.37 $Y2=1.667
r81 12 17 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=4.37 $Y=1.45
+ $X2=4.37 $Y2=1.235
r82 10 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.35 $Y=0.69
+ $X2=4.35 $Y2=1.085
r83 5 25 23.572 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=3.995 $Y=1.885
+ $X2=3.995 $Y2=1.667
r84 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.995 $Y=1.885
+ $X2=3.995 $Y2=2.46
r85 1 24 23.572 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=3.92 $Y=1.45 $X2=3.92
+ $Y2=1.667
r86 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.92 $Y=1.45 $X2=3.92
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%B1 1 3 4 5 6 8 9 11 12 14 15 16 21
c57 12 0 1.88567e-19 $X=5.865 $Y=1.885
r58 19 21 36.15 $w=6e-07 $l=4.5e-07 $layer=POLY_cond $X=5.542 $Y=1.165 $X2=5.542
+ $Y2=1.615
r59 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.615 $X2=6
+ $Y2=1.615
r60 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.57
+ $Y=1.615 $X2=5.57 $Y2=1.615
r61 12 21 46.1454 $w=3e-07 $l=4.37652e-07 $layer=POLY_cond $X=5.865 $Y=1.885
+ $X2=5.542 $Y2=1.615
r62 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.865 $Y=1.885
+ $X2=5.865 $Y2=2.46
r63 9 21 46.1454 $w=3e-07 $l=3.27399e-07 $layer=POLY_cond $X=5.415 $Y=1.885
+ $X2=5.542 $Y2=1.615
r64 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.415 $Y=1.885
+ $X2=5.415 $Y2=2.46
r65 6 19 37.3534 $w=6e-07 $l=3.57539e-07 $layer=POLY_cond $X=5.22 $Y=1.09
+ $X2=5.542 $Y2=1.165
r66 6 8 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.22 $Y=1.09 $X2=5.22
+ $Y2=0.69
r67 4 19 36.0747 $w=1.5e-07 $l=3.97e-07 $layer=POLY_cond $X=5.145 $Y=1.165
+ $X2=5.542 $Y2=1.165
r68 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.145 $Y=1.165
+ $X2=4.865 $Y2=1.165
r69 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.79 $Y=1.09
+ $X2=4.865 $Y2=1.165
r70 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.79 $Y=1.09 $X2=4.79
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%A1 1 3 6 8 10 13 15 16 24
c54 1 0 5.37684e-20 $X=6.315 $Y=1.885
r55 24 25 7.06933 $w=3.75e-07 $l=5.5e-08 $layer=POLY_cond $X=6.765 $Y=1.667
+ $X2=6.82 $Y2=1.667
r56 22 24 40.488 $w=3.75e-07 $l=3.15e-07 $layer=POLY_cond $X=6.45 $Y=1.667
+ $X2=6.765 $Y2=1.667
r57 20 22 7.712 $w=3.75e-07 $l=6e-08 $layer=POLY_cond $X=6.39 $Y=1.667 $X2=6.45
+ $Y2=1.667
r58 19 20 9.64 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=6.315 $Y=1.667
+ $X2=6.39 $Y2=1.667
r59 15 16 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=6.45 $Y=1.615
+ $X2=6.96 $Y2=1.615
r60 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.615 $X2=6.45 $Y2=1.615
r61 11 25 24.2915 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.82 $Y=1.45
+ $X2=6.82 $Y2=1.667
r62 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.82 $Y=1.45
+ $X2=6.82 $Y2=0.69
r63 8 24 24.2915 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.765 $Y=1.885
+ $X2=6.765 $Y2=1.667
r64 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.765 $Y=1.885
+ $X2=6.765 $Y2=2.46
r65 4 20 24.2915 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.39 $Y=1.45
+ $X2=6.39 $Y2=1.667
r66 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.39 $Y=1.45 $X2=6.39
+ $Y2=0.69
r67 1 19 24.2915 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.315 $Y=1.885
+ $X2=6.315 $Y2=1.667
r68 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.315 $Y=1.885
+ $X2=6.315 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%A2 2 3 5 8 11 12 14 17 19 20 30
c49 30 0 7.29804e-20 $X=7.68 $Y=1.425
c50 8 0 1.83628e-19 $X=7.25 $Y=0.69
r51 29 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.665 $Y=1.425
+ $X2=7.68 $Y2=1.425
r52 27 29 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=7.41 $Y=1.425
+ $X2=7.665 $Y2=1.425
r53 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.41
+ $Y=1.425 $X2=7.41 $Y2=1.425
r54 25 27 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=7.25 $Y=1.425
+ $X2=7.41 $Y2=1.425
r55 23 25 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.215 $Y=1.425
+ $X2=7.25 $Y2=1.425
r56 19 20 11.0407 $w=5.18e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.52
+ $X2=7.92 $Y2=1.52
r57 19 28 0.690045 $w=5.18e-07 $l=3e-08 $layer=LI1_cond $X=7.44 $Y=1.52 $X2=7.41
+ $Y2=1.52
r58 15 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.68 $Y=1.26
+ $X2=7.68 $Y2=1.425
r59 15 17 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=7.68 $Y=1.26
+ $X2=7.68 $Y2=0.69
r60 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.665 $Y=1.885
+ $X2=7.665 $Y2=2.46
r61 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.665 $Y=1.795
+ $X2=7.665 $Y2=1.885
r62 10 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.665 $Y=1.59
+ $X2=7.665 $Y2=1.425
r63 10 11 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=7.665 $Y=1.59
+ $X2=7.665 $Y2=1.795
r64 6 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.25 $Y=1.26
+ $X2=7.25 $Y2=1.425
r65 6 8 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=7.25 $Y=1.26 $X2=7.25
+ $Y2=0.69
r66 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.215 $Y=1.885
+ $X2=7.215 $Y2=2.46
r67 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.215 $Y=1.795 $X2=7.215
+ $Y2=1.885
r68 1 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.215 $Y=1.59
+ $X2=7.215 $Y2=1.425
r69 1 2 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=7.215 $Y=1.59
+ $X2=7.215 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%VPWR 1 2 3 4 5 18 22 26 32 36 39 40 42 43
+ 45 46 47 59 66 73 74 77 80
c101 32 0 1.88567e-19 $X=6.54 $Y=2.4
r102 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r103 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r104 74 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r105 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 71 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.525 $Y=3.33
+ $X2=7.4 $Y2=3.33
r107 71 73 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.525 $Y=3.33
+ $X2=7.92 $Y2=3.33
r108 70 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r109 70 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r111 67 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.54 $Y2=3.33
r112 67 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.96 $Y2=3.33
r113 66 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.275 $Y=3.33
+ $X2=7.4 $Y2=3.33
r114 66 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.275 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 65 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r116 64 65 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r117 61 64 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=6
+ $Y2=3.33
r118 61 62 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 59 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=3.33
+ $X2=6.54 $Y2=3.33
r120 59 64 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.375 $Y=3.33
+ $X2=6 $Y2=3.33
r121 58 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r123 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r124 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r127 47 65 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r128 47 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 45 57 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.39 $Y2=3.33
r131 44 61 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.64 $Y2=3.33
r132 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.39 $Y2=3.33
r133 42 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.45 $Y2=3.33
r135 41 57 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.45 $Y2=3.33
r137 39 50 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.24 $Y2=3.33
r138 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.51 $Y2=3.33
r139 38 54 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.51 $Y2=3.33
r141 34 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.4 $Y2=3.33
r142 34 36 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.4 $Y2=2.455
r143 30 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.54 $Y=3.245
+ $X2=6.54 $Y2=3.33
r144 30 32 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=6.54 $Y=3.245
+ $X2=6.54 $Y2=2.4
r145 26 29 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.39 $Y=1.985
+ $X2=2.39 $Y2=2.815
r146 24 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=3.245
+ $X2=2.39 $Y2=3.33
r147 24 29 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.39 $Y=3.245
+ $X2=2.39 $Y2=2.815
r148 20 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=3.245
+ $X2=1.45 $Y2=3.33
r149 20 22 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.45 $Y=3.245
+ $X2=1.45 $Y2=2.305
r150 16 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.51 $Y=3.245
+ $X2=0.51 $Y2=3.33
r151 16 18 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=0.51 $Y=3.245
+ $X2=0.51 $Y2=2.305
r152 5 36 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=7.29
+ $Y=1.96 $X2=7.44 $Y2=2.455
r153 4 32 300 $w=1.7e-07 $l=5.0951e-07 $layer=licon1_PDIFF $count=2 $X=6.39
+ $Y=1.96 $X2=6.54 $Y2=2.4
r154 3 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=1.84 $X2=2.35 $Y2=2.815
r155 3 26 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=1.84 $X2=2.35 $Y2=1.985
r156 2 22 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.3
+ $Y=1.84 $X2=1.45 $Y2=2.305
r157 1 18 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.425
+ $Y=1.84 $X2=0.55 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 39 43
+ 44 45 46
r78 45 46 8.42951 $w=5.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.387 $Y=1.295
+ $X2=0.387 $Y2=1.665
r79 42 46 3.07563 $w=5.23e-07 $l=1.35e-07 $layer=LI1_cond $X=0.387 $Y=1.8
+ $X2=0.387 $Y2=1.665
r80 41 45 3.7591 $w=5.23e-07 $l=1.65e-07 $layer=LI1_cond $X=0.387 $Y=1.13
+ $X2=0.387 $Y2=1.295
r81 37 39 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.32 $Y=0.96
+ $X2=2.32 $Y2=0.515
r82 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.9 $Y=1.985 $X2=1.9
+ $Y2=2.815
r83 31 33 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.9 $Y=1.97 $X2=1.9
+ $Y2=1.985
r84 30 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=1.045
+ $X2=1.54 $Y2=1.045
r85 29 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.195 $Y=1.045
+ $X2=2.32 $Y2=0.96
r86 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.195 $Y=1.045
+ $X2=1.665 $Y2=1.045
r87 25 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.96
+ $X2=1.54 $Y2=1.045
r88 25 27 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.54 $Y=0.96
+ $X2=1.54 $Y2=0.515
r89 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=1.885 $X2=1
+ $Y2=1.885
r90 23 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.735 $Y=1.885
+ $X2=1.9 $Y2=1.97
r91 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.735 $Y=1.885
+ $X2=1.165 $Y2=1.885
r92 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1 $Y=1.985 $X2=1
+ $Y2=2.815
r93 17 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1 $Y=1.97 $X2=1
+ $Y2=1.885
r94 17 19 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1 $Y=1.97 $X2=1
+ $Y2=1.985
r95 16 42 9.43933 $w=1.7e-07 $l=3.02529e-07 $layer=LI1_cond $X=0.65 $Y=1.885
+ $X2=0.387 $Y2=1.8
r96 15 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=1.885 $X2=1
+ $Y2=1.885
r97 15 16 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=1.885
+ $X2=0.65 $Y2=1.885
r98 14 41 9.43933 $w=1.7e-07 $l=3.02529e-07 $layer=LI1_cond $X=0.65 $Y=1.045
+ $X2=0.387 $Y2=1.13
r99 13 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=1.045
+ $X2=1.54 $Y2=1.045
r100 13 14 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.415 $Y=1.045
+ $X2=0.65 $Y2=1.045
r101 4 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=1.84 $X2=1.9 $Y2=2.815
r102 4 33 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=1.84 $X2=1.9 $Y2=1.985
r103 3 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.85
+ $Y=1.84 $X2=1 $Y2=2.815
r104 3 19 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.85
+ $Y=1.84 $X2=1 $Y2=1.985
r105 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.22
+ $Y=0.37 $X2=2.36 $Y2=0.515
r106 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.36
+ $Y=0.37 $X2=1.5 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%A_549_392# 1 2 3 12 14 15 18 22 26 28
r48 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.67 $Y=2.905
+ $X2=4.67 $Y2=2.455
r49 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.935 $Y=2.99
+ $X2=3.77 $Y2=2.99
r50 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.505 $Y=2.99
+ $X2=4.67 $Y2=2.905
r51 22 23 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.505 $Y=2.99
+ $X2=3.935 $Y2=2.99
r52 18 21 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=3.77 $Y=2.115 $X2=3.77
+ $Y2=2.815
r53 16 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=2.905
+ $X2=3.77 $Y2=2.99
r54 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.77 $Y=2.905 $X2=3.77
+ $Y2=2.815
r55 14 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=2.99
+ $X2=3.77 $Y2=2.99
r56 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.605 $Y=2.99
+ $X2=3.035 $Y2=2.99
r57 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.87 $Y=2.905
+ $X2=3.035 $Y2=2.99
r58 10 12 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.87 $Y=2.905
+ $X2=2.87 $Y2=2.455
r59 3 26 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=4.52
+ $Y=1.96 $X2=4.67 $Y2=2.455
r60 2 21 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.62
+ $Y=1.96 $X2=3.77 $Y2=2.815
r61 2 18 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=3.62
+ $Y=1.96 $X2=3.77 $Y2=2.115
r62 1 12 300 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.96 $X2=2.87 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%A_814_392# 1 2 9 14 16
c30 16 0 5.37684e-20 $X=5.64 $Y=2.115
r31 10 14 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=2.035
+ $X2=4.22 $Y2=2.035
r32 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.475 $Y=2.035
+ $X2=5.64 $Y2=2.035
r33 9 10 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=5.475 $Y=2.035
+ $X2=4.305 $Y2=2.035
r34 2 16 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=5.49
+ $Y=1.96 $X2=5.64 $Y2=2.115
r35 1 14 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=4.07
+ $Y=1.96 $X2=4.22 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%A_1013_392# 1 2 3 4 15 17 18 19 22 23 27 29
+ 31 33 38
r58 31 40 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=2.12 $X2=7.89
+ $Y2=2.035
r59 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.89 $Y=2.12
+ $X2=7.89 $Y2=2.815
r60 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=2.035
+ $X2=6.99 $Y2=2.035
r61 29 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.725 $Y=2.035
+ $X2=7.89 $Y2=2.035
r62 29 30 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.725 $Y=2.035
+ $X2=7.075 $Y2=2.035
r63 25 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=2.12 $X2=6.99
+ $Y2=2.035
r64 25 27 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.99 $Y=2.12
+ $X2=6.99 $Y2=2.815
r65 24 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=2.035
+ $X2=6.09 $Y2=2.035
r66 23 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=2.035
+ $X2=6.99 $Y2=2.035
r67 23 24 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.905 $Y=2.035
+ $X2=6.175 $Y2=2.035
r68 20 22 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.09 $Y=2.905 $X2=6.09
+ $Y2=2.815
r69 19 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=2.12 $X2=6.09
+ $Y2=2.035
r70 19 22 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.09 $Y=2.12
+ $X2=6.09 $Y2=2.815
r71 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.005 $Y=2.99
+ $X2=6.09 $Y2=2.905
r72 17 18 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.005 $Y=2.99
+ $X2=5.305 $Y2=2.99
r73 13 18 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=5.165 $Y=2.905
+ $X2=5.305 $Y2=2.99
r74 13 15 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=5.165 $Y=2.905
+ $X2=5.165 $Y2=2.455
r75 4 40 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=7.74
+ $Y=1.96 $X2=7.89 $Y2=2.115
r76 4 33 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=7.74
+ $Y=1.96 $X2=7.89 $Y2=2.815
r77 3 38 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.96 $X2=6.99 $Y2=2.115
r78 3 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.96 $X2=6.99 $Y2=2.815
r79 2 36 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.94
+ $Y=1.96 $X2=6.09 $Y2=2.115
r80 2 22 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.94
+ $Y=1.96 $X2=6.09 $Y2=2.815
r81 1 15 300 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=2 $X=5.065
+ $Y=1.96 $X2=5.19 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%VGND 1 2 3 4 5 6 7 24 28 30 34 36 40 44 48
+ 52 55 56 57 58 59 68 73 78 85 86 89 92 95 98 101
r114 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r115 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r116 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r117 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r118 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r119 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r120 86 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r121 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r122 83 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.63 $Y=0
+ $X2=7.465 $Y2=0
r123 83 85 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.63 $Y=0 $X2=7.92
+ $Y2=0
r124 82 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r125 82 99 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.52 $Y2=0
r126 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r127 79 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.6 $Y=0 $X2=5.435
+ $Y2=0
r128 79 81 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=5.6 $Y=0 $X2=6.96
+ $Y2=0
r129 78 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=7.465
+ $Y2=0
r130 78 81 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=6.96
+ $Y2=0
r131 77 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r132 77 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r133 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r134 74 95 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.57
+ $Y2=0
r135 74 76 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=5.04
+ $Y2=0
r136 73 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=0 $X2=5.435
+ $Y2=0
r137 73 76 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.27 $Y=0 $X2=5.04
+ $Y2=0
r138 69 92 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=3.7
+ $Y2=0
r139 69 71 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=4.08
+ $Y2=0
r140 68 95 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.4 $Y=0 $X2=4.57
+ $Y2=0
r141 68 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=0 $X2=4.08
+ $Y2=0
r142 67 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r143 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r144 63 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r145 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r146 59 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r147 59 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r148 59 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r149 57 66 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0
+ $X2=1.68 $Y2=0
r150 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=0 $X2=1.93
+ $Y2=0
r151 55 62 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r152 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r153 54 66 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=1.68 $Y2=0
r154 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r155 50 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.465 $Y=0.085
+ $X2=7.465 $Y2=0
r156 50 52 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=7.465 $Y=0.085
+ $X2=7.465 $Y2=0.585
r157 46 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=0.085
+ $X2=5.435 $Y2=0
r158 46 48 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.435 $Y=0.085
+ $X2=5.435 $Y2=0.515
r159 42 95 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=0.085
+ $X2=4.57 $Y2=0
r160 42 44 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=4.57 $Y=0.085
+ $X2=4.57 $Y2=0.495
r161 38 92 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0
r162 38 40 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.55
r163 37 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.75
+ $Y2=0
r164 36 92 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.53 $Y=0 $X2=3.7
+ $Y2=0
r165 36 37 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.53 $Y=0
+ $X2=2.875 $Y2=0
r166 32 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=0.085
+ $X2=2.75 $Y2=0
r167 32 34 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.75 $Y=0.085
+ $X2=2.75 $Y2=0.515
r168 31 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=0 $X2=1.93
+ $Y2=0
r169 30 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.75
+ $Y2=0
r170 30 31 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.625 $Y=0
+ $X2=2.015 $Y2=0
r171 26 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0
r172 26 28 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0.625
r173 22 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r174 22 24 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.625
r175 7 52 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=7.325
+ $Y=0.37 $X2=7.465 $Y2=0.585
r176 6 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.37 $X2=5.435 $Y2=0.515
r177 5 44 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.425
+ $Y=0.37 $X2=4.57 $Y2=0.495
r178 4 40 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=3.555
+ $Y=0.37 $X2=3.7 $Y2=0.55
r179 3 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.65
+ $Y=0.37 $X2=2.79 $Y2=0.515
r180 2 28 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.79
+ $Y=0.37 $X2=1.93 $Y2=0.625
r181 1 24 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=0.925
+ $Y=0.37 $X2=1.07 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_HS__A2111O_4%A_1210_74# 1 2 3 12 14 15 20 21 24
r36 22 24 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=7.935 $Y=0.92
+ $X2=7.935 $Y2=0.515
r37 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.81 $Y=1.005
+ $X2=7.935 $Y2=0.92
r38 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.81 $Y=1.005
+ $X2=7.12 $Y2=1.005
r39 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.035 $Y=0.92
+ $X2=7.12 $Y2=1.005
r40 17 19 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.035 $Y=0.92
+ $X2=7.035 $Y2=0.515
r41 16 19 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=7.035 $Y=0.455
+ $X2=7.035 $Y2=0.515
r42 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.95 $Y=0.37
+ $X2=7.035 $Y2=0.455
r43 14 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.95 $Y=0.37
+ $X2=6.34 $Y2=0.37
r44 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.175 $Y=0.455
+ $X2=6.34 $Y2=0.37
r45 10 12 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=6.175 $Y=0.455
+ $X2=6.175 $Y2=0.515
r46 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.755
+ $Y=0.37 $X2=7.895 $Y2=0.515
r47 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.895
+ $Y=0.37 $X2=7.035 $Y2=0.515
r48 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.05
+ $Y=0.37 $X2=6.175 $Y2=0.515
.ends

