* File: sky130_fd_sc_hs__dlxtn_4.pxi.spice
* Created: Tue Sep  1 20:03:09 2020
* 
x_PM_SKY130_FD_SC_HS__DLXTN_4%D N_D_M1011_g N_D_c_157_n N_D_c_161_n N_D_M1004_g
+ D N_D_c_158_n N_D_c_159_n PM_SKY130_FD_SC_HS__DLXTN_4%D
x_PM_SKY130_FD_SC_HS__DLXTN_4%GATE_N N_GATE_N_c_186_n N_GATE_N_M1019_g
+ N_GATE_N_M1017_g GATE_N PM_SKY130_FD_SC_HS__DLXTN_4%GATE_N
x_PM_SKY130_FD_SC_HS__DLXTN_4%A_230_424# N_A_230_424#_M1017_d
+ N_A_230_424#_M1019_d N_A_230_424#_c_236_n N_A_230_424#_M1006_g
+ N_A_230_424#_c_224_n N_A_230_424#_M1007_g N_A_230_424#_c_225_n
+ N_A_230_424#_M1001_g N_A_230_424#_c_226_n N_A_230_424#_c_237_n
+ N_A_230_424#_c_238_n N_A_230_424#_M1008_g N_A_230_424#_c_227_n
+ N_A_230_424#_c_228_n N_A_230_424#_c_229_n N_A_230_424#_c_230_n
+ N_A_230_424#_c_239_n N_A_230_424#_c_293_p N_A_230_424#_c_240_n
+ N_A_230_424#_c_241_n N_A_230_424#_c_242_n N_A_230_424#_c_243_n
+ N_A_230_424#_c_244_n N_A_230_424#_c_231_n N_A_230_424#_c_232_n
+ N_A_230_424#_c_233_n N_A_230_424#_c_234_n N_A_230_424#_c_235_n
+ PM_SKY130_FD_SC_HS__DLXTN_4%A_230_424#
x_PM_SKY130_FD_SC_HS__DLXTN_4%A_27_115# N_A_27_115#_M1011_s N_A_27_115#_M1004_s
+ N_A_27_115#_c_378_n N_A_27_115#_c_389_n N_A_27_115#_M1014_g
+ N_A_27_115#_c_379_n N_A_27_115#_M1002_g N_A_27_115#_c_390_n
+ N_A_27_115#_c_380_n N_A_27_115#_c_409_n N_A_27_115#_c_381_n
+ N_A_27_115#_c_382_n N_A_27_115#_c_383_n N_A_27_115#_c_384_n
+ N_A_27_115#_c_385_n N_A_27_115#_c_392_n N_A_27_115#_c_386_n
+ N_A_27_115#_c_387_n PM_SKY130_FD_SC_HS__DLXTN_4%A_27_115#
x_PM_SKY130_FD_SC_HS__DLXTN_4%A_369_392# N_A_369_392#_M1007_s
+ N_A_369_392#_M1006_s N_A_369_392#_c_493_n N_A_369_392#_M1018_g
+ N_A_369_392#_c_494_n N_A_369_392#_M1010_g N_A_369_392#_c_495_n
+ N_A_369_392#_c_502_n N_A_369_392#_c_496_n N_A_369_392#_c_497_n
+ N_A_369_392#_c_503_n N_A_369_392#_c_498_n N_A_369_392#_c_499_n
+ N_A_369_392#_c_500_n PM_SKY130_FD_SC_HS__DLXTN_4%A_369_392#
x_PM_SKY130_FD_SC_HS__DLXTN_4%A_840_395# N_A_840_395#_M1009_s
+ N_A_840_395#_M1012_d N_A_840_395#_c_601_n N_A_840_395#_M1020_g
+ N_A_840_395#_M1005_g N_A_840_395#_M1013_g N_A_840_395#_c_603_n
+ N_A_840_395#_M1000_g N_A_840_395#_c_591_n N_A_840_395#_M1016_g
+ N_A_840_395#_c_604_n N_A_840_395#_M1003_g N_A_840_395#_M1023_g
+ N_A_840_395#_c_605_n N_A_840_395#_M1021_g N_A_840_395#_M1025_g
+ N_A_840_395#_c_606_n N_A_840_395#_M1022_g N_A_840_395#_c_607_n
+ N_A_840_395#_c_595_n N_A_840_395#_c_596_n N_A_840_395#_c_608_n
+ N_A_840_395#_c_597_n N_A_840_395#_c_598_n N_A_840_395#_c_610_n
+ N_A_840_395#_c_599_n N_A_840_395#_c_650_p N_A_840_395#_c_600_n
+ PM_SKY130_FD_SC_HS__DLXTN_4%A_840_395#
x_PM_SKY130_FD_SC_HS__DLXTN_4%A_675_392# N_A_675_392#_M1001_d
+ N_A_675_392#_M1018_d N_A_675_392#_c_752_n N_A_675_392#_c_753_n
+ N_A_675_392#_M1012_g N_A_675_392#_M1009_g N_A_675_392#_M1024_g
+ N_A_675_392#_c_754_n N_A_675_392#_c_755_n N_A_675_392#_M1015_g
+ N_A_675_392#_c_745_n N_A_675_392#_c_746_n N_A_675_392#_c_747_n
+ N_A_675_392#_c_748_n N_A_675_392#_c_749_n N_A_675_392#_c_756_n
+ N_A_675_392#_c_750_n N_A_675_392#_c_751_n
+ PM_SKY130_FD_SC_HS__DLXTN_4%A_675_392#
x_PM_SKY130_FD_SC_HS__DLXTN_4%VPWR N_VPWR_M1004_d N_VPWR_M1006_d N_VPWR_M1020_d
+ N_VPWR_M1015_s N_VPWR_M1003_d N_VPWR_M1022_d N_VPWR_c_853_n N_VPWR_c_854_n
+ N_VPWR_c_855_n N_VPWR_c_856_n N_VPWR_c_857_n N_VPWR_c_858_n VPWR
+ N_VPWR_c_859_n N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n N_VPWR_c_863_n
+ N_VPWR_c_864_n N_VPWR_c_865_n N_VPWR_c_866_n N_VPWR_c_867_n N_VPWR_c_868_n
+ N_VPWR_c_869_n N_VPWR_c_852_n PM_SKY130_FD_SC_HS__DLXTN_4%VPWR
x_PM_SKY130_FD_SC_HS__DLXTN_4%Q N_Q_M1013_d N_Q_M1023_d N_Q_M1000_s N_Q_M1021_s
+ N_Q_c_954_n N_Q_c_961_n N_Q_c_962_n N_Q_c_955_n N_Q_c_956_n N_Q_c_957_n
+ N_Q_c_963_n N_Q_c_958_n N_Q_c_959_n Q Q Q N_Q_c_966_n
+ PM_SKY130_FD_SC_HS__DLXTN_4%Q
x_PM_SKY130_FD_SC_HS__DLXTN_4%VGND N_VGND_M1011_d N_VGND_M1007_d N_VGND_M1005_d
+ N_VGND_M1024_d N_VGND_M1016_s N_VGND_M1025_s N_VGND_c_1027_n N_VGND_c_1028_n
+ N_VGND_c_1029_n N_VGND_c_1030_n N_VGND_c_1031_n N_VGND_c_1032_n
+ N_VGND_c_1033_n N_VGND_c_1034_n N_VGND_c_1035_n VGND N_VGND_c_1036_n
+ N_VGND_c_1037_n N_VGND_c_1038_n N_VGND_c_1039_n N_VGND_c_1040_n
+ N_VGND_c_1041_n N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n
+ N_VGND_c_1045_n PM_SKY130_FD_SC_HS__DLXTN_4%VGND
cc_1 VNB N_D_M1011_g 0.0301791f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.85
cc_2 VNB N_D_c_157_n 0.00201979f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.955
cc_3 VNB N_D_c_158_n 0.00385705f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_D_c_159_n 0.060667f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.465
cc_5 VNB N_GATE_N_c_186_n 0.0147514f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_6 VNB N_GATE_N_M1017_g 0.0248735f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.955
cc_7 VNB GATE_N 0.00210952f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_8 VNB N_A_230_424#_c_224_n 0.0184509f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A_230_424#_c_225_n 0.0146603f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_10 VNB N_A_230_424#_c_226_n 0.010741f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.465
cc_11 VNB N_A_230_424#_c_227_n 0.0315798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_230_424#_c_228_n 0.0078699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_230_424#_c_229_n 0.00995015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_230_424#_c_230_n 0.00246166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_230_424#_c_231_n 0.0390372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_230_424#_c_232_n 5.47787e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_230_424#_c_233_n 0.00385597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_230_424#_c_234_n 0.0373933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_230_424#_c_235_n 0.0699059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_115#_c_378_n 0.00682663f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_21 VNB N_A_27_115#_c_379_n 0.0158604f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_22 VNB N_A_27_115#_c_380_n 0.00858581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_115#_c_381_n 0.0302799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_115#_c_382_n 0.00508052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_115#_c_383_n 0.023918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_115#_c_384_n 0.00292455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_115#_c_385_n 0.00224314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_115#_c_386_n 0.00833773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_115#_c_387_n 0.0611553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_369_392#_c_493_n 0.0210772f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.045
cc_31 VNB N_A_369_392#_c_494_n 0.0203856f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_A_369_392#_c_495_n 4.52811e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_369_392#_c_496_n 0.00222566f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_34 VNB N_A_369_392#_c_497_n 0.00678992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_369_392#_c_498_n 0.00365986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_369_392#_c_499_n 0.00796467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_369_392#_c_500_n 0.0480288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_840_395#_M1005_g 0.0448479f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_39 VNB N_A_840_395#_M1013_g 0.0247252f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_40 VNB N_A_840_395#_c_591_n 0.0248873f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_41 VNB N_A_840_395#_M1016_g 0.0223921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_840_395#_M1023_g 0.0217972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_840_395#_M1025_g 0.0243109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_840_395#_c_595_n 0.00214537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_840_395#_c_596_n 0.00197273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_840_395#_c_597_n 0.0121816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_840_395#_c_598_n 0.0105365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_840_395#_c_599_n 0.00409951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_840_395#_c_600_n 0.0679719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_675_392#_M1009_g 0.0272194f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_51 VNB N_A_675_392#_M1024_g 0.0240565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_675_392#_c_745_n 0.0071265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_675_392#_c_746_n 2.95717e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_675_392#_c_747_n 0.0027358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_675_392#_c_748_n 0.00356499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_675_392#_c_749_n 0.00933825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_675_392#_c_750_n 0.00418601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_675_392#_c_751_n 0.0430459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VPWR_c_852_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_Q_c_954_n 0.00299103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Q_c_955_n 0.00315465f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_62 VNB N_Q_c_956_n 0.00244574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_Q_c_957_n 0.00253236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_Q_c_958_n 0.00875216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_Q_c_959_n 0.00219521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB Q 0.0258426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1027_n 0.0163672f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_68 VNB N_VGND_c_1028_n 0.00988336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1029_n 0.0147111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1030_n 0.0061968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1031_n 0.00333063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1032_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1033_n 0.0296685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1034_n 0.0175031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1035_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1036_n 0.0195521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1037_n 0.0440818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1038_n 0.0436262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1039_n 0.0194943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1040_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1041_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1042_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1043_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1044_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1045_n 0.453881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VPB N_D_c_157_n 0.0236108f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.955
cc_87 VPB N_D_c_161_n 0.0269575f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.045
cc_88 VPB N_D_c_158_n 0.00761464f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_89 VPB N_GATE_N_c_186_n 0.0515183f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_90 VPB GATE_N 0.002419f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.54
cc_91 VPB N_A_230_424#_c_236_n 0.018527f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.045
cc_92 VPB N_A_230_424#_c_237_n 0.0367381f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_93 VPB N_A_230_424#_c_238_n 0.0209569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_230_424#_c_239_n 0.00668467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_230_424#_c_240_n 0.00564075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_230_424#_c_241_n 0.00210552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_230_424#_c_242_n 0.00750579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_230_424#_c_243_n 0.030543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_230_424#_c_244_n 0.00694013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_230_424#_c_232_n 0.00367977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_230_424#_c_233_n 0.00174569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_230_424#_c_234_n 0.0181944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_230_424#_c_235_n 0.0371045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_115#_c_378_n 0.00748721f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.54
cc_105 VPB N_A_27_115#_c_389_n 0.0229257f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.54
cc_106 VPB N_A_27_115#_c_390_n 0.0360197f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.465
cc_107 VPB N_A_27_115#_c_380_n 0.00559717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_115#_c_392_n 0.0156571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_369_392#_c_493_n 0.0340043f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.045
cc_110 VPB N_A_369_392#_c_502_n 0.0208346f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.465
cc_111 VPB N_A_369_392#_c_503_n 0.0071863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_369_392#_c_498_n 0.00263684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_840_395#_c_601_n 0.103121f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.045
cc_114 VPB N_A_840_395#_M1005_g 0.00568598f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_115 VPB N_A_840_395#_c_603_n 0.0169305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_840_395#_c_604_n 0.0154782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_840_395#_c_605_n 0.0148819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_840_395#_c_606_n 0.017188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_840_395#_c_607_n 0.00525346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_840_395#_c_608_n 0.00171897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_840_395#_c_597_n 0.00779621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_840_395#_c_610_n 0.0105894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_840_395#_c_600_n 0.0197739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_675_392#_c_752_n 0.0124334f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.54
cc_125 VPB N_A_675_392#_c_753_n 0.022635f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.54
cc_126 VPB N_A_675_392#_c_754_n 0.010912f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.665
cc_127 VPB N_A_675_392#_c_755_n 0.0229452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_675_392#_c_756_n 0.00162764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_675_392#_c_750_n 0.00325463f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_675_392#_c_751_n 0.0089239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_853_n 0.00970163f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.665
cc_132 VPB N_VPWR_c_854_n 0.0142812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_855_n 0.00841492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_856_n 0.00274039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_857_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_858_n 0.0341745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_859_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_860_n 0.0402815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_861_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_862_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_863_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_864_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_865_n 0.00864213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_866_n 0.0377908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_867_n 0.026624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_868_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_869_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_852_n 0.0868098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_Q_c_961_n 0.00226181f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.465
cc_150 VPB N_Q_c_962_n 0.00326984f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_151 VPB N_Q_c_963_n 0.00233217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB Q 0.00860207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB Q 0.0172459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_Q_c_966_n 0.00219771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 N_D_c_161_n N_GATE_N_c_186_n 0.0227883f $X=0.525 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_156 N_D_c_159_n N_GATE_N_c_186_n 0.0148841f $X=0.525 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_157 N_D_M1011_g N_GATE_N_M1017_g 0.0187327f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_158 N_D_c_159_n N_GATE_N_M1017_g 0.00470907f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_159 N_D_c_161_n N_A_230_424#_c_243_n 6.81629e-19 $X=0.525 $Y=2.045 $X2=0
+ $Y2=0
cc_160 N_D_c_161_n N_A_27_115#_c_390_n 0.0137802f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_161 N_D_M1011_g N_A_27_115#_c_380_n 0.00436712f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_162 N_D_c_158_n N_A_27_115#_c_380_n 0.036032f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_163 N_D_c_159_n N_A_27_115#_c_380_n 0.00955881f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_164 N_D_M1011_g N_A_27_115#_c_381_n 0.0278868f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_165 N_D_c_158_n N_A_27_115#_c_381_n 0.0279826f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_166 N_D_c_159_n N_A_27_115#_c_381_n 0.00435879f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_167 N_D_M1011_g N_A_27_115#_c_382_n 7.68306e-19 $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_168 N_D_c_157_n N_A_27_115#_c_392_n 0.00736553f $X=0.525 $Y=1.955 $X2=0 $Y2=0
cc_169 N_D_c_161_n N_A_27_115#_c_392_n 0.0140847f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_170 N_D_c_158_n N_A_27_115#_c_392_n 0.0260287f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_171 N_D_c_159_n N_A_27_115#_c_392_n 0.00146215f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_172 N_D_c_161_n N_VPWR_c_853_n 0.00737447f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_173 N_D_c_161_n N_VPWR_c_859_n 0.00445602f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_174 N_D_c_161_n N_VPWR_c_852_n 0.00861384f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_175 N_D_M1011_g N_VGND_c_1027_n 0.00130869f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_176 N_D_M1011_g N_VGND_c_1036_n 0.00341528f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_177 N_D_M1011_g N_VGND_c_1045_n 0.0048347f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_178 N_GATE_N_c_186_n N_A_230_424#_c_228_n 0.00354352f $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_179 N_GATE_N_M1017_g N_A_230_424#_c_228_n 0.00566256f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_180 GATE_N N_A_230_424#_c_228_n 0.0141427f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_181 N_GATE_N_M1017_g N_A_230_424#_c_229_n 0.00371584f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_182 N_GATE_N_c_186_n N_A_230_424#_c_230_n 0.00135088f $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_183 N_GATE_N_M1017_g N_A_230_424#_c_230_n 0.00359662f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_184 GATE_N N_A_230_424#_c_230_n 0.0260997f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_185 N_GATE_N_c_186_n N_A_230_424#_c_239_n 2.30203e-19 $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_186 N_GATE_N_c_186_n N_A_230_424#_c_243_n 0.0188904f $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_187 GATE_N N_A_230_424#_c_243_n 0.0106287f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_188 N_GATE_N_c_186_n N_A_230_424#_c_244_n 0.00795499f $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_189 N_GATE_N_M1017_g N_A_230_424#_c_231_n 0.0155068f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_190 N_GATE_N_c_186_n N_A_230_424#_c_235_n 0.0149176f $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_191 GATE_N N_A_230_424#_c_235_n 2.97788e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_192 N_GATE_N_c_186_n N_A_27_115#_c_390_n 6.6422e-19 $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_193 N_GATE_N_c_186_n N_A_27_115#_c_380_n 0.00370557f $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_194 N_GATE_N_M1017_g N_A_27_115#_c_380_n 0.00516253f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_195 GATE_N N_A_27_115#_c_380_n 0.022773f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_196 N_GATE_N_M1017_g N_A_27_115#_c_409_n 0.0140794f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_197 GATE_N N_A_27_115#_c_409_n 0.00313461f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_198 N_GATE_N_M1017_g N_A_27_115#_c_381_n 0.00639387f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_199 N_GATE_N_M1017_g N_A_27_115#_c_382_n 0.00773574f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_200 N_GATE_N_c_186_n N_A_27_115#_c_392_n 0.00425246f $X=1.075 $Y=2.045 $X2=0
+ $Y2=0
cc_201 N_GATE_N_c_186_n N_VPWR_c_853_n 0.00737447f $X=1.075 $Y=2.045 $X2=0 $Y2=0
cc_202 N_GATE_N_c_186_n N_VPWR_c_860_n 0.00445602f $X=1.075 $Y=2.045 $X2=0 $Y2=0
cc_203 N_GATE_N_c_186_n N_VPWR_c_852_n 0.00862626f $X=1.075 $Y=2.045 $X2=0 $Y2=0
cc_204 N_GATE_N_M1017_g N_VGND_c_1027_n 5.5317e-19 $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_205 N_GATE_N_M1017_g N_VGND_c_1037_n 0.00318127f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_206 N_GATE_N_M1017_g N_VGND_c_1045_n 0.00438121f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_207 N_A_230_424#_c_235_n N_A_27_115#_c_378_n 0.008372f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_208 N_A_230_424#_c_236_n N_A_27_115#_c_389_n 0.0242388f $X=2.215 $Y=1.885
+ $X2=0 $Y2=0
cc_209 N_A_230_424#_c_239_n N_A_27_115#_c_389_n 0.0136166f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_210 N_A_230_424#_c_241_n N_A_27_115#_c_389_n 0.00118311f $X=3.16 $Y=2.99
+ $X2=0 $Y2=0
cc_211 N_A_230_424#_c_224_n N_A_27_115#_c_379_n 0.00442933f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_212 N_A_230_424#_c_225_n N_A_27_115#_c_379_n 0.0227686f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_213 N_A_230_424#_c_243_n N_A_27_115#_c_390_n 0.00419773f $X=1.3 $Y=2.265
+ $X2=0 $Y2=0
cc_214 N_A_230_424#_c_228_n N_A_27_115#_c_380_n 0.00915345f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_215 N_A_230_424#_M1017_d N_A_27_115#_c_409_n 0.00613024f $X=1.16 $Y=0.57
+ $X2=0 $Y2=0
cc_216 N_A_230_424#_c_228_n N_A_27_115#_c_409_n 0.00997713f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_217 N_A_230_424#_c_229_n N_A_27_115#_c_409_n 0.00618319f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_218 N_A_230_424#_c_231_n N_A_27_115#_c_409_n 2.54774e-19 $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_219 N_A_230_424#_c_228_n N_A_27_115#_c_381_n 0.00659465f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_220 N_A_230_424#_M1017_d N_A_27_115#_c_382_n 0.00339584f $X=1.16 $Y=0.57
+ $X2=0 $Y2=0
cc_221 N_A_230_424#_c_224_n N_A_27_115#_c_383_n 0.0157054f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_222 N_A_230_424#_c_228_n N_A_27_115#_c_383_n 0.00552911f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_223 N_A_230_424#_c_229_n N_A_27_115#_c_383_n 0.0169889f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_224 N_A_230_424#_c_231_n N_A_27_115#_c_383_n 0.00199179f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_225 N_A_230_424#_c_224_n N_A_27_115#_c_385_n 0.00730669f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_226 N_A_230_424#_c_243_n N_A_27_115#_c_392_n 9.83506e-19 $X=1.3 $Y=2.265
+ $X2=0 $Y2=0
cc_227 N_A_230_424#_c_235_n N_A_27_115#_c_386_n 0.00293022f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_228 N_A_230_424#_c_224_n N_A_27_115#_c_387_n 0.00242956f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_229 N_A_230_424#_c_227_n N_A_27_115#_c_387_n 0.0227686f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_230 N_A_230_424#_c_235_n N_A_27_115#_c_387_n 0.0131368f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_231 N_A_230_424#_c_239_n N_A_369_392#_M1006_s 0.00788967f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_232 N_A_230_424#_c_237_n N_A_369_392#_c_493_n 0.012f $X=3.87 $Y=2.375 $X2=0
+ $Y2=0
cc_233 N_A_230_424#_c_238_n N_A_369_392#_c_493_n 0.0124548f $X=3.87 $Y=2.465
+ $X2=0 $Y2=0
cc_234 N_A_230_424#_c_227_n N_A_369_392#_c_493_n 6.79409e-19 $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_235 N_A_230_424#_c_239_n N_A_369_392#_c_493_n 0.00142562f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_236 N_A_230_424#_c_293_p N_A_369_392#_c_493_n 0.0052118f $X=3.075 $Y=2.905
+ $X2=0 $Y2=0
cc_237 N_A_230_424#_c_240_n N_A_369_392#_c_493_n 0.0134991f $X=4.05 $Y=2.99
+ $X2=0 $Y2=0
cc_238 N_A_230_424#_c_234_n N_A_369_392#_c_493_n 0.0173938f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_239 N_A_230_424#_c_225_n N_A_369_392#_c_494_n 0.00527673f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_240 N_A_230_424#_c_227_n N_A_369_392#_c_494_n 0.00161375f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_241 N_A_230_424#_c_233_n N_A_369_392#_c_494_n 2.45027e-19 $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_242 N_A_230_424#_c_234_n N_A_369_392#_c_494_n 0.00312708f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_243 N_A_230_424#_c_224_n N_A_369_392#_c_495_n 0.00940637f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_244 N_A_230_424#_c_229_n N_A_369_392#_c_495_n 0.044954f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_245 N_A_230_424#_c_230_n N_A_369_392#_c_495_n 0.0289818f $X=1.685 $Y=1.57
+ $X2=0 $Y2=0
cc_246 N_A_230_424#_c_231_n N_A_369_392#_c_495_n 0.00156461f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_247 N_A_230_424#_c_235_n N_A_369_392#_c_495_n 0.0278331f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_248 N_A_230_424#_c_239_n N_A_369_392#_c_502_n 0.0263218f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_249 N_A_230_424#_c_235_n N_A_369_392#_c_502_n 0.00411697f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_250 N_A_230_424#_c_225_n N_A_369_392#_c_497_n 0.0173976f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_251 N_A_230_424#_c_227_n N_A_369_392#_c_497_n 6.03378e-19 $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_252 N_A_230_424#_c_236_n N_A_369_392#_c_503_n 0.0129511f $X=2.215 $Y=1.885
+ $X2=0 $Y2=0
cc_253 N_A_230_424#_c_239_n N_A_369_392#_c_503_n 0.0285858f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_254 N_A_230_424#_c_244_n N_A_369_392#_c_503_n 0.0311123f $X=1.395 $Y=2.1
+ $X2=0 $Y2=0
cc_255 N_A_230_424#_c_232_n N_A_369_392#_c_503_n 0.00896259f $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_256 N_A_230_424#_c_235_n N_A_369_392#_c_503_n 0.0183834f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_257 N_A_230_424#_c_237_n N_A_369_392#_c_498_n 2.90563e-19 $X=3.87 $Y=2.375
+ $X2=0 $Y2=0
cc_258 N_A_230_424#_c_234_n N_A_369_392#_c_498_n 3.62762e-19 $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_259 N_A_230_424#_c_225_n N_A_369_392#_c_499_n 0.00376963f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_260 N_A_230_424#_c_226_n N_A_369_392#_c_499_n 0.00118688f $X=3.855 $Y=1.405
+ $X2=0 $Y2=0
cc_261 N_A_230_424#_c_225_n N_A_369_392#_c_500_n 0.00586767f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_262 N_A_230_424#_c_237_n N_A_840_395#_c_601_n 0.026732f $X=3.87 $Y=2.375
+ $X2=0 $Y2=0
cc_263 N_A_230_424#_c_238_n N_A_840_395#_c_601_n 0.0272633f $X=3.87 $Y=2.465
+ $X2=0 $Y2=0
cc_264 N_A_230_424#_c_240_n N_A_840_395#_c_601_n 0.00351728f $X=4.05 $Y=2.99
+ $X2=0 $Y2=0
cc_265 N_A_230_424#_c_242_n N_A_840_395#_c_601_n 0.0301913f $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_266 N_A_230_424#_c_233_n N_A_840_395#_c_601_n 0.0012023f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_267 N_A_230_424#_c_234_n N_A_840_395#_c_601_n 0.0101586f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_268 N_A_230_424#_c_242_n N_A_840_395#_M1005_g 6.0243e-19 $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_269 N_A_230_424#_c_233_n N_A_840_395#_M1005_g 7.74691e-19 $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_270 N_A_230_424#_c_234_n N_A_840_395#_M1005_g 0.0136936f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_271 N_A_230_424#_c_242_n N_A_840_395#_c_607_n 0.0249855f $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_272 N_A_230_424#_c_240_n N_A_675_392#_M1018_d 0.00343217f $X=4.05 $Y=2.99
+ $X2=0 $Y2=0
cc_273 N_A_230_424#_c_227_n N_A_675_392#_c_745_n 0.00249179f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_274 N_A_230_424#_c_233_n N_A_675_392#_c_745_n 0.0154026f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_275 N_A_230_424#_c_234_n N_A_675_392#_c_745_n 0.00598369f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_276 N_A_230_424#_c_225_n N_A_675_392#_c_746_n 0.00514497f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_277 N_A_230_424#_c_227_n N_A_675_392#_c_746_n 0.00126393f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_278 N_A_230_424#_c_227_n N_A_675_392#_c_747_n 0.00254147f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_279 N_A_230_424#_c_226_n N_A_675_392#_c_748_n 0.00128751f $X=3.855 $Y=1.405
+ $X2=0 $Y2=0
cc_280 N_A_230_424#_c_233_n N_A_675_392#_c_748_n 0.0206617f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_281 N_A_230_424#_c_234_n N_A_675_392#_c_748_n 0.00196022f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_282 N_A_230_424#_c_237_n N_A_675_392#_c_756_n 0.00987965f $X=3.87 $Y=2.375
+ $X2=0 $Y2=0
cc_283 N_A_230_424#_c_238_n N_A_675_392#_c_756_n 0.012397f $X=3.87 $Y=2.465
+ $X2=0 $Y2=0
cc_284 N_A_230_424#_c_239_n N_A_675_392#_c_756_n 0.0127867f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_285 N_A_230_424#_c_293_p N_A_675_392#_c_756_n 0.0117819f $X=3.075 $Y=2.905
+ $X2=0 $Y2=0
cc_286 N_A_230_424#_c_240_n N_A_675_392#_c_756_n 0.0302235f $X=4.05 $Y=2.99
+ $X2=0 $Y2=0
cc_287 N_A_230_424#_c_242_n N_A_675_392#_c_756_n 0.0494584f $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_288 N_A_230_424#_c_225_n N_A_675_392#_c_750_n 6.76373e-19 $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_289 N_A_230_424#_c_226_n N_A_675_392#_c_750_n 0.00615882f $X=3.855 $Y=1.405
+ $X2=0 $Y2=0
cc_290 N_A_230_424#_c_237_n N_A_675_392#_c_750_n 0.00755818f $X=3.87 $Y=2.375
+ $X2=0 $Y2=0
cc_291 N_A_230_424#_c_227_n N_A_675_392#_c_750_n 0.0117959f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_292 N_A_230_424#_c_233_n N_A_675_392#_c_750_n 0.0494584f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_293 N_A_230_424#_c_234_n N_A_675_392#_c_750_n 0.00971643f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_294 N_A_230_424#_c_239_n N_VPWR_M1006_d 0.0129815f $X=2.99 $Y=2.475 $X2=0
+ $Y2=0
cc_295 N_A_230_424#_c_243_n N_VPWR_c_853_n 0.0285454f $X=1.3 $Y=2.265 $X2=0
+ $Y2=0
cc_296 N_A_230_424#_c_236_n N_VPWR_c_854_n 0.00622405f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_297 N_A_230_424#_c_239_n N_VPWR_c_854_n 0.0316438f $X=2.99 $Y=2.475 $X2=0
+ $Y2=0
cc_298 N_A_230_424#_c_241_n N_VPWR_c_854_n 0.0120577f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_299 N_A_230_424#_c_236_n N_VPWR_c_860_n 0.00469064f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_300 N_A_230_424#_c_243_n N_VPWR_c_860_n 0.0230718f $X=1.3 $Y=2.265 $X2=0
+ $Y2=0
cc_301 N_A_230_424#_c_238_n N_VPWR_c_866_n 0.00278271f $X=3.87 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A_230_424#_c_240_n N_VPWR_c_866_n 0.0685372f $X=4.05 $Y=2.99 $X2=0
+ $Y2=0
cc_303 N_A_230_424#_c_241_n N_VPWR_c_866_n 0.0121935f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_304 N_A_230_424#_c_240_n N_VPWR_c_867_n 0.0125323f $X=4.05 $Y=2.99 $X2=0
+ $Y2=0
cc_305 N_A_230_424#_c_236_n N_VPWR_c_852_n 0.0049649f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_306 N_A_230_424#_c_238_n N_VPWR_c_852_n 0.00354684f $X=3.87 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_230_424#_c_239_n N_VPWR_c_852_n 0.0323484f $X=2.99 $Y=2.475 $X2=0
+ $Y2=0
cc_308 N_A_230_424#_c_240_n N_VPWR_c_852_n 0.0386705f $X=4.05 $Y=2.99 $X2=0
+ $Y2=0
cc_309 N_A_230_424#_c_241_n N_VPWR_c_852_n 0.00661049f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_310 N_A_230_424#_c_243_n N_VPWR_c_852_n 0.0190639f $X=1.3 $Y=2.265 $X2=0
+ $Y2=0
cc_311 N_A_230_424#_c_239_n A_591_392# 0.00457165f $X=2.99 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_312 N_A_230_424#_c_293_p A_591_392# 0.00389072f $X=3.075 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_313 N_A_230_424#_c_240_n A_591_392# 2.67089e-19 $X=4.05 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_314 N_A_230_424#_c_240_n A_789_508# 0.00179331f $X=4.05 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A_230_424#_c_242_n A_789_508# 0.00349116f $X=4.135 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_316 N_A_230_424#_c_224_n N_VGND_c_1028_n 0.00195643f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_317 N_A_230_424#_c_225_n N_VGND_c_1028_n 3.35588e-19 $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_318 N_A_230_424#_c_224_n N_VGND_c_1037_n 0.00278271f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_319 N_A_230_424#_c_225_n N_VGND_c_1038_n 9.44495e-19 $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_320 N_A_230_424#_c_224_n N_VGND_c_1045_n 0.00363426f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_321 N_A_27_115#_c_383_n N_A_369_392#_M1007_s 0.00441657f $X=2.475 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_322 N_A_27_115#_c_378_n N_A_369_392#_c_493_n 0.018592f $X=2.88 $Y=1.795 $X2=0
+ $Y2=0
cc_323 N_A_27_115#_c_389_n N_A_369_392#_c_493_n 0.0524617f $X=2.88 $Y=1.885
+ $X2=0 $Y2=0
cc_324 N_A_27_115#_c_386_n N_A_369_392#_c_493_n 2.74972e-19 $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_325 N_A_27_115#_c_387_n N_A_369_392#_c_493_n 0.0104126f $X=2.88 $Y=1.33 $X2=0
+ $Y2=0
cc_326 N_A_27_115#_c_378_n N_A_369_392#_c_495_n 9.39281e-19 $X=2.88 $Y=1.795
+ $X2=0 $Y2=0
cc_327 N_A_27_115#_c_383_n N_A_369_392#_c_495_n 0.0144209f $X=2.475 $Y=0.34
+ $X2=0 $Y2=0
cc_328 N_A_27_115#_c_385_n N_A_369_392#_c_495_n 0.0265397f $X=2.56 $Y=1.22 $X2=0
+ $Y2=0
cc_329 N_A_27_115#_c_386_n N_A_369_392#_c_495_n 0.0265613f $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_330 N_A_27_115#_c_387_n N_A_369_392#_c_495_n 2.87669e-19 $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_331 N_A_27_115#_c_378_n N_A_369_392#_c_502_n 0.00571054f $X=2.88 $Y=1.795
+ $X2=0 $Y2=0
cc_332 N_A_27_115#_c_389_n N_A_369_392#_c_502_n 0.00817455f $X=2.88 $Y=1.885
+ $X2=0 $Y2=0
cc_333 N_A_27_115#_c_386_n N_A_369_392#_c_502_n 0.0395884f $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_334 N_A_27_115#_c_387_n N_A_369_392#_c_502_n 0.00785784f $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_335 N_A_27_115#_c_379_n N_A_369_392#_c_496_n 0.00147103f $X=3.215 $Y=1.11
+ $X2=0 $Y2=0
cc_336 N_A_27_115#_c_389_n N_A_369_392#_c_503_n 0.00157273f $X=2.88 $Y=1.885
+ $X2=0 $Y2=0
cc_337 N_A_27_115#_c_378_n N_A_369_392#_c_498_n 0.00122989f $X=2.88 $Y=1.795
+ $X2=0 $Y2=0
cc_338 N_A_27_115#_c_386_n N_A_369_392#_c_498_n 0.00521207f $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_339 N_A_27_115#_c_387_n N_A_369_392#_c_498_n 7.06729e-19 $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_340 N_A_27_115#_c_379_n N_A_369_392#_c_499_n 0.00497566f $X=3.215 $Y=1.11
+ $X2=0 $Y2=0
cc_341 N_A_27_115#_c_385_n N_A_369_392#_c_499_n 0.00474149f $X=2.56 $Y=1.22
+ $X2=0 $Y2=0
cc_342 N_A_27_115#_c_386_n N_A_369_392#_c_499_n 0.0122394f $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_343 N_A_27_115#_c_387_n N_A_369_392#_c_499_n 0.00129573f $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_344 N_A_27_115#_c_389_n N_A_675_392#_c_756_n 0.00176562f $X=2.88 $Y=1.885
+ $X2=0 $Y2=0
cc_345 N_A_27_115#_c_390_n N_VPWR_c_853_n 0.0266809f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_346 N_A_27_115#_c_392_n N_VPWR_c_853_n 0.0121673f $X=0.71 $Y=2.035 $X2=0
+ $Y2=0
cc_347 N_A_27_115#_c_389_n N_VPWR_c_854_n 0.0108748f $X=2.88 $Y=1.885 $X2=0
+ $Y2=0
cc_348 N_A_27_115#_c_390_n N_VPWR_c_859_n 0.0145938f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_349 N_A_27_115#_c_389_n N_VPWR_c_866_n 0.00413917f $X=2.88 $Y=1.885 $X2=0
+ $Y2=0
cc_350 N_A_27_115#_c_389_n N_VPWR_c_852_n 0.00398447f $X=2.88 $Y=1.885 $X2=0
+ $Y2=0
cc_351 N_A_27_115#_c_390_n N_VPWR_c_852_n 0.0120466f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_352 N_A_27_115#_c_380_n N_VGND_M1011_d 0.00236148f $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_353 N_A_27_115#_c_409_n N_VGND_M1011_d 0.007918f $X=1.145 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_354 N_A_27_115#_c_381_n N_VGND_M1011_d 0.00690665f $X=0.795 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_355 N_A_27_115#_c_383_n N_VGND_M1007_d 6.47853e-19 $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_356 N_A_27_115#_c_385_n N_VGND_M1007_d 0.0110808f $X=2.56 $Y=1.22 $X2=0 $Y2=0
cc_357 N_A_27_115#_c_409_n N_VGND_c_1027_n 0.0121815f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_358 N_A_27_115#_c_381_n N_VGND_c_1027_n 0.0143324f $X=0.795 $Y=0.745 $X2=0
+ $Y2=0
cc_359 N_A_27_115#_c_382_n N_VGND_c_1027_n 0.0045384f $X=1.23 $Y=0.66 $X2=0
+ $Y2=0
cc_360 N_A_27_115#_c_384_n N_VGND_c_1027_n 0.0139003f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_361 N_A_27_115#_c_379_n N_VGND_c_1028_n 0.0092719f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_362 N_A_27_115#_c_383_n N_VGND_c_1028_n 0.0148948f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_363 N_A_27_115#_c_385_n N_VGND_c_1028_n 0.0477502f $X=2.56 $Y=1.22 $X2=0
+ $Y2=0
cc_364 N_A_27_115#_c_386_n N_VGND_c_1028_n 0.0155155f $X=2.835 $Y=1.385 $X2=0
+ $Y2=0
cc_365 N_A_27_115#_c_387_n N_VGND_c_1028_n 0.00987931f $X=2.88 $Y=1.33 $X2=0
+ $Y2=0
cc_366 N_A_27_115#_c_381_n N_VGND_c_1036_n 0.0103718f $X=0.795 $Y=0.745 $X2=0
+ $Y2=0
cc_367 N_A_27_115#_c_409_n N_VGND_c_1037_n 0.00257035f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_368 N_A_27_115#_c_383_n N_VGND_c_1037_n 0.086417f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_369 N_A_27_115#_c_384_n N_VGND_c_1037_n 0.0120335f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_370 N_A_27_115#_c_379_n N_VGND_c_1038_n 0.00539704f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_371 N_A_27_115#_c_379_n N_VGND_c_1045_n 0.0052351f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_372 N_A_27_115#_c_409_n N_VGND_c_1045_n 0.00589268f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_373 N_A_27_115#_c_381_n N_VGND_c_1045_n 0.0164998f $X=0.795 $Y=0.745 $X2=0
+ $Y2=0
cc_374 N_A_27_115#_c_383_n N_VGND_c_1045_n 0.049532f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_375 N_A_27_115#_c_384_n N_VGND_c_1045_n 0.00658039f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_376 N_A_369_392#_c_500_n N_A_840_395#_M1005_g 0.0424929f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_377 N_A_369_392#_c_497_n N_A_675_392#_M1001_d 0.00252704f $X=4.28 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_378 N_A_369_392#_c_500_n N_A_675_392#_M1009_g 0.00207621f $X=4.4 $Y=0.34
+ $X2=0 $Y2=0
cc_379 N_A_369_392#_c_494_n N_A_675_392#_c_745_n 0.0151004f $X=4.4 $Y=0.505
+ $X2=0 $Y2=0
cc_380 N_A_369_392#_c_497_n N_A_675_392#_c_745_n 0.0316369f $X=4.28 $Y=0.34
+ $X2=0 $Y2=0
cc_381 N_A_369_392#_c_500_n N_A_675_392#_c_745_n 0.00447421f $X=4.4 $Y=0.34
+ $X2=0 $Y2=0
cc_382 N_A_369_392#_c_497_n N_A_675_392#_c_746_n 0.0105171f $X=4.28 $Y=0.34
+ $X2=0 $Y2=0
cc_383 N_A_369_392#_c_499_n N_A_675_392#_c_746_n 0.0146188f $X=3.375 $Y=1.47
+ $X2=0 $Y2=0
cc_384 N_A_369_392#_c_494_n N_A_675_392#_c_747_n 0.0012686f $X=4.4 $Y=0.505
+ $X2=0 $Y2=0
cc_385 N_A_369_392#_c_493_n N_A_675_392#_c_756_n 0.010685f $X=3.3 $Y=1.885 $X2=0
+ $Y2=0
cc_386 N_A_369_392#_c_498_n N_A_675_392#_c_756_n 0.0134669f $X=3.375 $Y=1.635
+ $X2=0 $Y2=0
cc_387 N_A_369_392#_c_493_n N_A_675_392#_c_750_n 0.00502278f $X=3.3 $Y=1.885
+ $X2=0 $Y2=0
cc_388 N_A_369_392#_c_494_n N_A_675_392#_c_750_n 6.66919e-19 $X=4.4 $Y=0.505
+ $X2=0 $Y2=0
cc_389 N_A_369_392#_c_498_n N_A_675_392#_c_750_n 0.031936f $X=3.375 $Y=1.635
+ $X2=0 $Y2=0
cc_390 N_A_369_392#_c_499_n N_A_675_392#_c_750_n 0.0250348f $X=3.375 $Y=1.47
+ $X2=0 $Y2=0
cc_391 N_A_369_392#_c_493_n N_VPWR_c_854_n 2.61619e-19 $X=3.3 $Y=1.885 $X2=0
+ $Y2=0
cc_392 N_A_369_392#_c_493_n N_VPWR_c_866_n 0.00278271f $X=3.3 $Y=1.885 $X2=0
+ $Y2=0
cc_393 N_A_369_392#_c_493_n N_VPWR_c_852_n 0.00354684f $X=3.3 $Y=1.885 $X2=0
+ $Y2=0
cc_394 N_A_369_392#_c_502_n N_VGND_c_1028_n 0.00457271f $X=3.21 $Y=1.805 $X2=0
+ $Y2=0
cc_395 N_A_369_392#_c_496_n N_VGND_c_1028_n 0.0159466f $X=3.485 $Y=0.38 $X2=0
+ $Y2=0
cc_396 N_A_369_392#_c_499_n N_VGND_c_1028_n 0.0209764f $X=3.375 $Y=1.47 $X2=0
+ $Y2=0
cc_397 N_A_369_392#_c_497_n N_VGND_c_1029_n 0.0098708f $X=4.28 $Y=0.34 $X2=0
+ $Y2=0
cc_398 N_A_369_392#_c_500_n N_VGND_c_1029_n 0.00431935f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_399 N_A_369_392#_c_496_n N_VGND_c_1038_n 0.0121867f $X=3.485 $Y=0.38 $X2=0
+ $Y2=0
cc_400 N_A_369_392#_c_497_n N_VGND_c_1038_n 0.062486f $X=4.28 $Y=0.34 $X2=0
+ $Y2=0
cc_401 N_A_369_392#_c_500_n N_VGND_c_1038_n 0.00730902f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_402 N_A_369_392#_c_496_n N_VGND_c_1045_n 0.00660921f $X=3.485 $Y=0.38 $X2=0
+ $Y2=0
cc_403 N_A_369_392#_c_497_n N_VGND_c_1045_n 0.0348893f $X=4.28 $Y=0.34 $X2=0
+ $Y2=0
cc_404 N_A_369_392#_c_500_n N_VGND_c_1045_n 0.0113113f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_405 N_A_369_392#_c_499_n A_658_79# 0.00247748f $X=3.375 $Y=1.47 $X2=-0.19
+ $Y2=-0.245
cc_406 N_A_840_395#_c_601_n N_A_675_392#_c_752_n 0.0108689f $X=4.29 $Y=2.465
+ $X2=0 $Y2=0
cc_407 N_A_840_395#_c_610_n N_A_675_392#_c_752_n 0.00501737f $X=5.48 $Y=2.265
+ $X2=0 $Y2=0
cc_408 N_A_840_395#_c_601_n N_A_675_392#_c_753_n 0.00796086f $X=4.29 $Y=2.465
+ $X2=0 $Y2=0
cc_409 N_A_840_395#_c_607_n N_A_675_392#_c_753_n 0.0226192f $X=5.315 $Y=2.14
+ $X2=0 $Y2=0
cc_410 N_A_840_395#_c_610_n N_A_675_392#_c_753_n 0.00106588f $X=5.48 $Y=2.265
+ $X2=0 $Y2=0
cc_411 N_A_840_395#_M1005_g N_A_675_392#_M1009_g 0.0178603f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_412 N_A_840_395#_c_595_n N_A_675_392#_M1009_g 0.00687953f $X=5.485 $Y=0.54
+ $X2=0 $Y2=0
cc_413 N_A_840_395#_c_596_n N_A_675_392#_M1009_g 9.92594e-19 $X=5.745 $Y=1.32
+ $X2=0 $Y2=0
cc_414 N_A_840_395#_c_599_n N_A_675_392#_M1009_g 0.00431125f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_415 N_A_840_395#_M1013_g N_A_675_392#_M1024_g 0.0239087f $X=6.215 $Y=0.74
+ $X2=0 $Y2=0
cc_416 N_A_840_395#_c_596_n N_A_675_392#_M1024_g 0.00552835f $X=5.745 $Y=1.32
+ $X2=0 $Y2=0
cc_417 N_A_840_395#_c_599_n N_A_675_392#_M1024_g 0.0120291f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_418 N_A_840_395#_c_603_n N_A_675_392#_c_754_n 0.00907633f $X=6.23 $Y=1.765
+ $X2=0 $Y2=0
cc_419 N_A_840_395#_c_608_n N_A_675_392#_c_754_n 0.00255388f $X=5.745 $Y=1.82
+ $X2=0 $Y2=0
cc_420 N_A_840_395#_c_610_n N_A_675_392#_c_754_n 0.00517991f $X=5.48 $Y=2.265
+ $X2=0 $Y2=0
cc_421 N_A_840_395#_c_603_n N_A_675_392#_c_755_n 0.0083341f $X=6.23 $Y=1.765
+ $X2=0 $Y2=0
cc_422 N_A_840_395#_c_610_n N_A_675_392#_c_755_n 0.0143589f $X=5.48 $Y=2.265
+ $X2=0 $Y2=0
cc_423 N_A_840_395#_M1005_g N_A_675_392#_c_745_n 0.00733517f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_424 N_A_840_395#_M1005_g N_A_675_392#_c_747_n 0.00826027f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_425 N_A_840_395#_c_599_n N_A_675_392#_c_747_n 0.00244264f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_426 N_A_840_395#_c_601_n N_A_675_392#_c_748_n 0.0034639f $X=4.29 $Y=2.465
+ $X2=0 $Y2=0
cc_427 N_A_840_395#_M1005_g N_A_675_392#_c_748_n 0.00512512f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_428 N_A_840_395#_c_607_n N_A_675_392#_c_748_n 0.00868744f $X=5.315 $Y=2.14
+ $X2=0 $Y2=0
cc_429 N_A_840_395#_M1005_g N_A_675_392#_c_749_n 0.0152674f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_430 N_A_840_395#_c_607_n N_A_675_392#_c_749_n 0.0294526f $X=5.315 $Y=2.14
+ $X2=0 $Y2=0
cc_431 N_A_840_395#_c_610_n N_A_675_392#_c_749_n 0.01476f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_432 N_A_840_395#_c_599_n N_A_675_392#_c_749_n 0.0126845f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_433 N_A_840_395#_c_650_p N_A_675_392#_c_749_n 0.0277655f $X=5.745 $Y=1.485
+ $X2=0 $Y2=0
cc_434 N_A_840_395#_c_601_n N_A_675_392#_c_756_n 2.35511e-19 $X=4.29 $Y=2.465
+ $X2=0 $Y2=0
cc_435 N_A_840_395#_c_601_n N_A_675_392#_c_750_n 4.15014e-19 $X=4.29 $Y=2.465
+ $X2=0 $Y2=0
cc_436 N_A_840_395#_M1005_g N_A_675_392#_c_751_n 0.0186005f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_437 N_A_840_395#_c_608_n N_A_675_392#_c_751_n 0.00389059f $X=5.745 $Y=1.82
+ $X2=0 $Y2=0
cc_438 N_A_840_395#_c_597_n N_A_675_392#_c_751_n 0.0150167f $X=6.305 $Y=1.485
+ $X2=0 $Y2=0
cc_439 N_A_840_395#_c_610_n N_A_675_392#_c_751_n 0.00393379f $X=5.48 $Y=2.265
+ $X2=0 $Y2=0
cc_440 N_A_840_395#_c_599_n N_A_675_392#_c_751_n 0.00257893f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_441 N_A_840_395#_c_650_p N_A_675_392#_c_751_n 0.0142276f $X=5.745 $Y=1.485
+ $X2=0 $Y2=0
cc_442 N_A_840_395#_c_607_n N_VPWR_M1020_d 0.00293121f $X=5.315 $Y=2.14 $X2=0
+ $Y2=0
cc_443 N_A_840_395#_c_603_n N_VPWR_c_855_n 0.00259104f $X=6.23 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_A_840_395#_c_598_n N_VPWR_c_855_n 0.0108616f $X=7.325 $Y=1.485 $X2=0
+ $Y2=0
cc_445 N_A_840_395#_c_610_n N_VPWR_c_855_n 0.00158095f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_446 N_A_840_395#_c_603_n N_VPWR_c_856_n 5.16951e-19 $X=6.23 $Y=1.765 $X2=0
+ $Y2=0
cc_447 N_A_840_395#_c_604_n N_VPWR_c_856_n 0.0141189f $X=6.755 $Y=1.765 $X2=0
+ $Y2=0
cc_448 N_A_840_395#_c_605_n N_VPWR_c_856_n 0.0138152f $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_449 N_A_840_395#_c_606_n N_VPWR_c_856_n 5.40442e-19 $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_450 N_A_840_395#_c_605_n N_VPWR_c_858_n 4.98648e-19 $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_451 N_A_840_395#_c_606_n N_VPWR_c_858_n 0.0116621f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_452 N_A_840_395#_c_610_n N_VPWR_c_861_n 0.0146357f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_453 N_A_840_395#_c_603_n N_VPWR_c_862_n 0.00461464f $X=6.23 $Y=1.765 $X2=0
+ $Y2=0
cc_454 N_A_840_395#_c_604_n N_VPWR_c_862_n 0.00413917f $X=6.755 $Y=1.765 $X2=0
+ $Y2=0
cc_455 N_A_840_395#_c_605_n N_VPWR_c_863_n 0.00413917f $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_456 N_A_840_395#_c_606_n N_VPWR_c_863_n 0.00413917f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_457 N_A_840_395#_c_601_n N_VPWR_c_866_n 0.00455353f $X=4.29 $Y=2.465 $X2=0
+ $Y2=0
cc_458 N_A_840_395#_c_601_n N_VPWR_c_867_n 0.0122177f $X=4.29 $Y=2.465 $X2=0
+ $Y2=0
cc_459 N_A_840_395#_c_607_n N_VPWR_c_867_n 0.0386877f $X=5.315 $Y=2.14 $X2=0
+ $Y2=0
cc_460 N_A_840_395#_c_610_n N_VPWR_c_867_n 0.0188056f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_461 N_A_840_395#_c_601_n N_VPWR_c_852_n 0.00929693f $X=4.29 $Y=2.465 $X2=0
+ $Y2=0
cc_462 N_A_840_395#_c_603_n N_VPWR_c_852_n 0.00908949f $X=6.23 $Y=1.765 $X2=0
+ $Y2=0
cc_463 N_A_840_395#_c_604_n N_VPWR_c_852_n 0.00818402f $X=6.755 $Y=1.765 $X2=0
+ $Y2=0
cc_464 N_A_840_395#_c_605_n N_VPWR_c_852_n 0.00817726f $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_465 N_A_840_395#_c_606_n N_VPWR_c_852_n 0.00817726f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_466 N_A_840_395#_c_610_n N_VPWR_c_852_n 0.0121141f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_467 N_A_840_395#_M1013_g N_Q_c_954_n 0.00944159f $X=6.215 $Y=0.74 $X2=0 $Y2=0
cc_468 N_A_840_395#_M1016_g N_Q_c_954_n 0.00350623f $X=6.735 $Y=0.74 $X2=0 $Y2=0
cc_469 N_A_840_395#_c_603_n N_Q_c_961_n 3.1841e-19 $X=6.23 $Y=1.765 $X2=0 $Y2=0
cc_470 N_A_840_395#_c_591_n N_Q_c_961_n 0.00807936f $X=6.66 $Y=1.485 $X2=0 $Y2=0
cc_471 N_A_840_395#_c_598_n N_Q_c_961_n 0.0277922f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_472 N_A_840_395#_c_610_n N_Q_c_961_n 0.00410663f $X=5.48 $Y=2.265 $X2=0 $Y2=0
cc_473 N_A_840_395#_c_603_n N_Q_c_962_n 4.83474e-19 $X=6.23 $Y=1.765 $X2=0 $Y2=0
cc_474 N_A_840_395#_c_604_n N_Q_c_962_n 0.00564841f $X=6.755 $Y=1.765 $X2=0
+ $Y2=0
cc_475 N_A_840_395#_M1016_g N_Q_c_955_n 0.0148325f $X=6.735 $Y=0.74 $X2=0 $Y2=0
cc_476 N_A_840_395#_M1023_g N_Q_c_955_n 0.0127761f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_477 N_A_840_395#_c_598_n N_Q_c_955_n 0.049875f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_478 N_A_840_395#_c_600_n N_Q_c_955_n 0.00224206f $X=7.64 $Y=1.542 $X2=0 $Y2=0
cc_479 N_A_840_395#_M1013_g N_Q_c_956_n 0.00366127f $X=6.215 $Y=0.74 $X2=0 $Y2=0
cc_480 N_A_840_395#_c_591_n N_Q_c_956_n 0.00442617f $X=6.66 $Y=1.485 $X2=0 $Y2=0
cc_481 N_A_840_395#_c_598_n N_Q_c_956_n 0.0293689f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_482 N_A_840_395#_c_599_n N_Q_c_956_n 0.00593633f $X=5.745 $Y=1.065 $X2=0
+ $Y2=0
cc_483 N_A_840_395#_M1023_g N_Q_c_957_n 4.44219e-19 $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_484 N_A_840_395#_M1025_g N_Q_c_957_n 4.74419e-19 $X=7.64 $Y=0.74 $X2=0 $Y2=0
cc_485 N_A_840_395#_c_605_n N_Q_c_963_n 3.85296e-19 $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_486 N_A_840_395#_c_606_n N_Q_c_963_n 3.85296e-19 $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_487 N_A_840_395#_M1025_g N_Q_c_958_n 0.0171357f $X=7.64 $Y=0.74 $X2=0 $Y2=0
cc_488 N_A_840_395#_c_600_n N_Q_c_958_n 7.24638e-19 $X=7.64 $Y=1.542 $X2=0 $Y2=0
cc_489 N_A_840_395#_c_598_n N_Q_c_959_n 0.016446f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_490 N_A_840_395#_c_600_n N_Q_c_959_n 0.00337787f $X=7.64 $Y=1.542 $X2=0 $Y2=0
cc_491 N_A_840_395#_M1025_g Q 0.0112315f $X=7.64 $Y=0.74 $X2=0 $Y2=0
cc_492 N_A_840_395#_c_606_n Q 0.00214581f $X=7.655 $Y=1.765 $X2=0 $Y2=0
cc_493 N_A_840_395#_c_598_n Q 0.0168437f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_494 N_A_840_395#_c_600_n Q 0.0105311f $X=7.64 $Y=1.542 $X2=0 $Y2=0
cc_495 N_A_840_395#_c_606_n Q 0.0223034f $X=7.655 $Y=1.765 $X2=0 $Y2=0
cc_496 N_A_840_395#_c_600_n Q 0.00105441f $X=7.64 $Y=1.542 $X2=0 $Y2=0
cc_497 N_A_840_395#_c_591_n N_Q_c_966_n 5.00849e-19 $X=6.66 $Y=1.485 $X2=0 $Y2=0
cc_498 N_A_840_395#_c_604_n N_Q_c_966_n 0.0150075f $X=6.755 $Y=1.765 $X2=0 $Y2=0
cc_499 N_A_840_395#_c_605_n N_Q_c_966_n 0.0129286f $X=7.205 $Y=1.765 $X2=0 $Y2=0
cc_500 N_A_840_395#_c_598_n N_Q_c_966_n 0.0629677f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_501 N_A_840_395#_c_600_n N_Q_c_966_n 0.0155978f $X=7.64 $Y=1.542 $X2=0 $Y2=0
cc_502 N_A_840_395#_M1005_g N_VGND_c_1029_n 0.00349542f $X=4.76 $Y=0.825 $X2=0
+ $Y2=0
cc_503 N_A_840_395#_c_595_n N_VGND_c_1029_n 0.0215088f $X=5.485 $Y=0.54 $X2=0
+ $Y2=0
cc_504 N_A_840_395#_c_599_n N_VGND_c_1029_n 0.00358005f $X=5.745 $Y=1.065 $X2=0
+ $Y2=0
cc_505 N_A_840_395#_M1013_g N_VGND_c_1030_n 0.00739063f $X=6.215 $Y=0.74 $X2=0
+ $Y2=0
cc_506 N_A_840_395#_c_595_n N_VGND_c_1030_n 0.0163189f $X=5.485 $Y=0.54 $X2=0
+ $Y2=0
cc_507 N_A_840_395#_c_598_n N_VGND_c_1030_n 0.00973029f $X=7.325 $Y=1.485 $X2=0
+ $Y2=0
cc_508 N_A_840_395#_c_599_n N_VGND_c_1030_n 0.00182821f $X=5.745 $Y=1.065 $X2=0
+ $Y2=0
cc_509 N_A_840_395#_M1013_g N_VGND_c_1031_n 6.65972e-19 $X=6.215 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_A_840_395#_M1016_g N_VGND_c_1031_n 0.0099317f $X=6.735 $Y=0.74 $X2=0
+ $Y2=0
cc_511 N_A_840_395#_M1023_g N_VGND_c_1031_n 0.00988667f $X=7.165 $Y=0.74 $X2=0
+ $Y2=0
cc_512 N_A_840_395#_M1025_g N_VGND_c_1031_n 4.5982e-19 $X=7.64 $Y=0.74 $X2=0
+ $Y2=0
cc_513 N_A_840_395#_M1025_g N_VGND_c_1033_n 0.00497413f $X=7.64 $Y=0.74 $X2=0
+ $Y2=0
cc_514 N_A_840_395#_c_595_n N_VGND_c_1034_n 0.00990263f $X=5.485 $Y=0.54 $X2=0
+ $Y2=0
cc_515 N_A_840_395#_M1005_g N_VGND_c_1038_n 0.00399533f $X=4.76 $Y=0.825 $X2=0
+ $Y2=0
cc_516 N_A_840_395#_M1013_g N_VGND_c_1039_n 0.00434272f $X=6.215 $Y=0.74 $X2=0
+ $Y2=0
cc_517 N_A_840_395#_M1016_g N_VGND_c_1039_n 0.00383152f $X=6.735 $Y=0.74 $X2=0
+ $Y2=0
cc_518 N_A_840_395#_M1023_g N_VGND_c_1040_n 0.00383152f $X=7.165 $Y=0.74 $X2=0
+ $Y2=0
cc_519 N_A_840_395#_M1025_g N_VGND_c_1040_n 0.00460063f $X=7.64 $Y=0.74 $X2=0
+ $Y2=0
cc_520 N_A_840_395#_M1005_g N_VGND_c_1045_n 0.00472204f $X=4.76 $Y=0.825 $X2=0
+ $Y2=0
cc_521 N_A_840_395#_M1013_g N_VGND_c_1045_n 0.00826226f $X=6.215 $Y=0.74 $X2=0
+ $Y2=0
cc_522 N_A_840_395#_M1016_g N_VGND_c_1045_n 0.00758371f $X=6.735 $Y=0.74 $X2=0
+ $Y2=0
cc_523 N_A_840_395#_M1023_g N_VGND_c_1045_n 0.00757973f $X=7.165 $Y=0.74 $X2=0
+ $Y2=0
cc_524 N_A_840_395#_M1025_g N_VGND_c_1045_n 0.00911274f $X=7.64 $Y=0.74 $X2=0
+ $Y2=0
cc_525 N_A_840_395#_c_595_n N_VGND_c_1045_n 0.0089622f $X=5.485 $Y=0.54 $X2=0
+ $Y2=0
cc_526 N_A_675_392#_c_755_n N_VPWR_c_855_n 0.00256351f $X=5.725 $Y=2.045 $X2=0
+ $Y2=0
cc_527 N_A_675_392#_c_753_n N_VPWR_c_861_n 0.00460063f $X=5.22 $Y=2.045 $X2=0
+ $Y2=0
cc_528 N_A_675_392#_c_755_n N_VPWR_c_861_n 0.00461464f $X=5.725 $Y=2.045 $X2=0
+ $Y2=0
cc_529 N_A_675_392#_c_753_n N_VPWR_c_867_n 0.00447129f $X=5.22 $Y=2.045 $X2=0
+ $Y2=0
cc_530 N_A_675_392#_c_755_n N_VPWR_c_867_n 3.36554e-19 $X=5.725 $Y=2.045 $X2=0
+ $Y2=0
cc_531 N_A_675_392#_c_753_n N_VPWR_c_852_n 0.0090472f $X=5.22 $Y=2.045 $X2=0
+ $Y2=0
cc_532 N_A_675_392#_c_755_n N_VPWR_c_852_n 0.00908891f $X=5.725 $Y=2.045 $X2=0
+ $Y2=0
cc_533 N_A_675_392#_M1024_g N_Q_c_954_n 9.40157e-19 $X=5.7 $Y=0.715 $X2=0 $Y2=0
cc_534 N_A_675_392#_M1009_g N_VGND_c_1029_n 0.00607982f $X=5.27 $Y=0.715 $X2=0
+ $Y2=0
cc_535 N_A_675_392#_c_745_n N_VGND_c_1029_n 0.0146621f $X=4.55 $Y=0.89 $X2=0
+ $Y2=0
cc_536 N_A_675_392#_c_749_n N_VGND_c_1029_n 0.0160858f $X=5.325 $Y=1.485 $X2=0
+ $Y2=0
cc_537 N_A_675_392#_M1009_g N_VGND_c_1030_n 4.73318e-19 $X=5.27 $Y=0.715 $X2=0
+ $Y2=0
cc_538 N_A_675_392#_M1024_g N_VGND_c_1030_n 0.00930995f $X=5.7 $Y=0.715 $X2=0
+ $Y2=0
cc_539 N_A_675_392#_M1009_g N_VGND_c_1034_n 0.00534051f $X=5.27 $Y=0.715 $X2=0
+ $Y2=0
cc_540 N_A_675_392#_M1024_g N_VGND_c_1034_n 0.00465077f $X=5.7 $Y=0.715 $X2=0
+ $Y2=0
cc_541 N_A_675_392#_c_745_n N_VGND_c_1038_n 0.00333424f $X=4.55 $Y=0.89 $X2=0
+ $Y2=0
cc_542 N_A_675_392#_M1009_g N_VGND_c_1045_n 0.00537853f $X=5.27 $Y=0.715 $X2=0
+ $Y2=0
cc_543 N_A_675_392#_M1024_g N_VGND_c_1045_n 0.00451796f $X=5.7 $Y=0.715 $X2=0
+ $Y2=0
cc_544 N_A_675_392#_c_745_n N_VGND_c_1045_n 0.00882318f $X=4.55 $Y=0.89 $X2=0
+ $Y2=0
cc_545 N_A_675_392#_c_745_n A_895_123# 0.00190356f $X=4.55 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_546 N_VPWR_c_855_n N_Q_c_962_n 0.00158095f $X=5.98 $Y=2.325 $X2=0 $Y2=0
cc_547 N_VPWR_c_856_n N_Q_c_962_n 0.0315588f $X=6.98 $Y=2.265 $X2=0 $Y2=0
cc_548 N_VPWR_c_862_n N_Q_c_962_n 0.0146357f $X=6.815 $Y=3.33 $X2=0 $Y2=0
cc_549 N_VPWR_c_852_n N_Q_c_962_n 0.0121141f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_550 N_VPWR_c_856_n N_Q_c_963_n 0.0315168f $X=6.98 $Y=2.265 $X2=0 $Y2=0
cc_551 N_VPWR_c_858_n N_Q_c_963_n 0.0255132f $X=7.88 $Y=2.405 $X2=0 $Y2=0
cc_552 N_VPWR_c_863_n N_Q_c_963_n 0.0101736f $X=7.715 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_852_n N_Q_c_963_n 0.0084208f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_554 N_VPWR_M1022_d Q 0.00454904f $X=7.73 $Y=1.84 $X2=0 $Y2=0
cc_555 N_VPWR_c_858_n Q 0.0221872f $X=7.88 $Y=2.405 $X2=0 $Y2=0
cc_556 N_VPWR_M1003_d N_Q_c_966_n 0.00197722f $X=6.83 $Y=1.84 $X2=0 $Y2=0
cc_557 N_VPWR_c_856_n N_Q_c_966_n 0.0171813f $X=6.98 $Y=2.265 $X2=0 $Y2=0
cc_558 N_Q_c_955_n N_VGND_M1016_s 0.00176461f $X=7.295 $Y=1.065 $X2=0 $Y2=0
cc_559 N_Q_c_958_n N_VGND_M1025_s 0.00371016f $X=7.805 $Y=1.065 $X2=0 $Y2=0
cc_560 N_Q_c_954_n N_VGND_c_1030_n 0.0336294f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_561 N_Q_c_954_n N_VGND_c_1031_n 0.0180579f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_562 N_Q_c_955_n N_VGND_c_1031_n 0.0170777f $X=7.295 $Y=1.065 $X2=0 $Y2=0
cc_563 N_Q_c_957_n N_VGND_c_1031_n 0.017215f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_564 N_Q_c_957_n N_VGND_c_1033_n 0.0175659f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_565 N_Q_c_958_n N_VGND_c_1033_n 0.0234209f $X=7.805 $Y=1.065 $X2=0 $Y2=0
cc_566 N_Q_c_954_n N_VGND_c_1039_n 0.0154563f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_567 N_Q_c_957_n N_VGND_c_1040_n 0.011066f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_568 N_Q_c_954_n N_VGND_c_1045_n 0.012737f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_569 N_Q_c_957_n N_VGND_c_1045_n 0.00915947f $X=7.38 $Y=0.515 $X2=0 $Y2=0
