* File: sky130_fd_sc_hs__ha_4.spice
* Created: Tue Sep  1 20:06:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__ha_4.pex.spice"
.subckt sky130_fd_sc_hs__ha_4  VNB VPB B A VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1016 N_A_27_125#_M1016_d N_A_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0912 PD=1.85 PS=0.925 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1021 N_A_27_125#_M1021_d N_A_M1021_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0912 PD=0.92 PS=0.925 NRD=0 NRS=0.936 M=1 R=4.26667 SA=75000.6
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_A_27_125#_M1021_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1004_d N_B_M1009_g N_A_27_125#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0992 PD=0.92 PS=0.95 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_294_392#_M1023_d N_A_435_99#_M1023_g N_A_27_125#_M1009_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1024 AS=0.0992 PD=0.96 PS=0.95 NRD=7.488 NRS=5.616 M=1
+ R=4.26667 SA=75002 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1025 N_A_294_392#_M1023_d N_A_435_99#_M1025_g N_A_27_125#_M1025_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1024 AS=0.2144 PD=0.96 PS=1.95 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75002.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1002 N_A_435_99#_M1002_d N_B_M1002_g N_A_707_119#_M1002_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1856 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1005 N_A_435_99#_M1002_d N_B_M1005_g N_A_707_119#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_707_119#_M1005_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.112 PD=0.99 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1006_d N_A_M1012_g N_A_707_119#_M1012_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.176 PD=0.99 PS=1.83 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_A_435_99#_M1010_g N_COUT_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2035 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_435_99#_M1013_g N_COUT_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75003 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1013_d N_A_435_99#_M1030_g N_COUT_M1030_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1033_d N_A_435_99#_M1033_g N_COUT_M1030_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1033_d N_A_294_392#_M1008_g N_SUM_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_A_294_392#_M1020_g N_SUM_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1020_d N_A_294_392#_M1024_g N_SUM_M1024_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.14985 PD=1.09 PS=1.145 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1028_d N_A_294_392#_M1028_g N_SUM_M1024_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.14985 PD=2.05 PS=1.145 NRD=0 NRS=8.916 M=1 R=4.93333
+ SA=75003.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_VPWR_M1026_d N_A_M1026_g N_A_27_392#_M1026_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.285 PD=1.3 PS=2.57 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1027 N_VPWR_M1026_d N_A_M1027_g N_A_27_392#_M1027_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.7
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1031 N_A_294_392#_M1031_d N_B_M1031_g N_A_27_392#_M1027_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1034 N_A_294_392#_M1031_d N_B_M1034_g N_A_27_392#_M1034_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.285 PD=1.3 PS=2.57 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1014 N_A_294_392#_M1014_d N_A_435_99#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.2394 PD=1.14 PS=2.25 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75005.6 A=0.126 P=1.98 MULT=1
MM1015 N_A_294_392#_M1014_d N_A_435_99#_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75000.7 SB=75005.1 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1015_s N_B_M1000_g N_A_435_99#_M1000_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.222537 PD=1.14 PS=1.58 NRD=2.3443 NRS=21.0987 M=1 R=5.6
+ SA=75001.1 SB=75004.7 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_B_M1018_g N_A_435_99#_M1000_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.222537 PD=1.14 PS=1.58 NRD=2.3443 NRS=49.2303 M=1 R=5.6
+ SA=75001.4 SB=75004.2 A=0.126 P=1.98 MULT=1
MM1003 N_A_435_99#_M1003_d N_A_M1003_g N_VPWR_M1018_d VPB PSHORT L=0.15 W=0.84
+ AD=0.175875 AS=0.126 PD=1.425 PS=1.14 NRD=36.1889 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75003.8 A=0.126 P=1.98 MULT=1
MM1011 N_A_435_99#_M1003_d N_A_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=0.84
+ AD=0.175875 AS=0.234 PD=1.425 PS=1.39714 NRD=0 NRS=52.4217 M=1 R=5.6
+ SA=75002.1 SB=75004.4 A=0.126 P=1.98 MULT=1
MM1017 N_COUT_M1017_d N_A_435_99#_M1017_g N_VPWR_M1011_s VPB PSHORT L=0.15
+ W=1.12 AD=0.2576 AS=0.312 PD=1.58 PS=1.86286 NRD=29.0181 NRS=13.1793 M=1
+ R=7.46667 SA=75002.1 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1022 N_COUT_M1017_d N_A_435_99#_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.15
+ W=1.12 AD=0.2576 AS=0.168 PD=1.58 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75002.7 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1029 N_COUT_M1029_d N_A_435_99#_M1029_g N_VPWR_M1022_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1032 N_COUT_M1029_d N_A_435_99#_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.6 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1032_s N_A_294_392#_M1001_g N_SUM_M1001_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.1 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A_294_392#_M1007_g N_SUM_M1001_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1007_d N_A_294_392#_M1019_g N_SUM_M1019_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3136 PD=1.42 PS=1.68 NRD=1.7533 NRS=28.1316 M=1 R=7.46667
+ SA=75005 SB=75000.9 A=0.168 P=2.54 MULT=1
MM1035 N_VPWR_M1035_d N_A_294_392#_M1035_g N_SUM_M1019_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.3136 PD=2.83 PS=1.68 NRD=1.7533 NRS=21.0987 M=1
+ R=7.46667 SA=75005.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX36_noxref VNB VPB NWDIODE A=19.5501 P=24.79
c_97 VNB 0 2.61855e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__ha_4.pxi.spice"
*
.ends
*
*
