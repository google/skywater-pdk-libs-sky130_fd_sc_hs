* File: sky130_fd_sc_hs__o211a_1.pxi.spice
* Created: Thu Aug 27 20:56:42 2020
* 
x_PM_SKY130_FD_SC_HS__O211A_1%A_83_264# N_A_83_264#_M1000_d N_A_83_264#_M1001_d
+ N_A_83_264#_M1009_d N_A_83_264#_M1008_g N_A_83_264#_c_70_n N_A_83_264#_M1005_g
+ N_A_83_264#_c_65_n N_A_83_264#_c_66_n N_A_83_264#_c_72_n N_A_83_264#_c_80_p
+ N_A_83_264#_c_128_p N_A_83_264#_c_73_n N_A_83_264#_c_67_n N_A_83_264#_c_97_p
+ N_A_83_264#_c_96_p N_A_83_264#_c_100_p N_A_83_264#_c_75_n N_A_83_264#_c_76_n
+ N_A_83_264#_c_124_p N_A_83_264#_c_68_n N_A_83_264#_c_77_n N_A_83_264#_c_69_n
+ PM_SKY130_FD_SC_HS__O211A_1%A_83_264#
x_PM_SKY130_FD_SC_HS__O211A_1%A1 N_A1_M1002_g N_A1_c_177_n N_A1_M1007_g A1
+ N_A1_c_175_n N_A1_c_176_n PM_SKY130_FD_SC_HS__O211A_1%A1
x_PM_SKY130_FD_SC_HS__O211A_1%A2 N_A2_c_212_n N_A2_c_213_n N_A2_c_218_n
+ N_A2_M1001_g N_A2_M1006_g A2 A2 A2 N_A2_c_216_n PM_SKY130_FD_SC_HS__O211A_1%A2
x_PM_SKY130_FD_SC_HS__O211A_1%B1 N_B1_c_255_n N_B1_M1003_g N_B1_M1004_g B1
+ N_B1_c_254_n PM_SKY130_FD_SC_HS__O211A_1%B1
x_PM_SKY130_FD_SC_HS__O211A_1%C1 N_C1_M1000_g N_C1_c_289_n N_C1_M1009_g C1
+ PM_SKY130_FD_SC_HS__O211A_1%C1
x_PM_SKY130_FD_SC_HS__O211A_1%X N_X_M1008_s N_X_M1005_s N_X_c_315_n N_X_c_316_n
+ X X X X N_X_c_317_n PM_SKY130_FD_SC_HS__O211A_1%X
x_PM_SKY130_FD_SC_HS__O211A_1%VPWR N_VPWR_M1005_d N_VPWR_M1003_d N_VPWR_c_342_n
+ VPWR N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_341_n N_VPWR_c_346_n
+ N_VPWR_c_347_n N_VPWR_c_348_n PM_SKY130_FD_SC_HS__O211A_1%VPWR
x_PM_SKY130_FD_SC_HS__O211A_1%VGND N_VGND_M1008_d N_VGND_M1002_d N_VGND_c_384_n
+ N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n VGND N_VGND_c_388_n
+ N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n PM_SKY130_FD_SC_HS__O211A_1%VGND
x_PM_SKY130_FD_SC_HS__O211A_1%A_257_136# N_A_257_136#_M1002_s
+ N_A_257_136#_M1006_d N_A_257_136#_c_423_n N_A_257_136#_c_427_n
+ N_A_257_136#_c_424_n N_A_257_136#_c_441_n N_A_257_136#_c_444_n
+ N_A_257_136#_c_432_n PM_SKY130_FD_SC_HS__O211A_1%A_257_136#
cc_1 VNB N_A_83_264#_M1008_g 0.0317094f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_83_264#_c_65_n 0.0169813f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.542
cc_3 VNB N_A_83_264#_c_66_n 0.00990888f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.65
cc_4 VNB N_A_83_264#_c_67_n 0.0050774f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=1.94
cc_5 VNB N_A_83_264#_c_68_n 0.0523754f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.485
cc_6 VNB N_A_83_264#_c_69_n 0.0317075f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.855
cc_7 VNB N_A1_M1002_g 0.0244149f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=1.96
cc_8 VNB N_A1_c_175_n 0.0353192f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_9 VNB N_A1_c_176_n 0.00479049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_c_212_n 0.00654074f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=0.68
cc_11 VNB N_A2_c_213_n 0.00879931f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=1.96
cc_12 VNB N_A2_M1006_g 0.014291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A2 0.0364706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_216_n 0.0503218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1004_g 0.0219731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB B1 0.00132948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_254_n 0.0305665f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_18 VNB N_C1_M1000_g 0.0268341f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=1.96
cc_19 VNB N_C1_c_289_n 0.0198909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB C1 0.0121714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_315_n 0.0265914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_316_n 0.0137581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_317_n 0.0249595f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=1.235
cc_24 VNB N_VPWR_c_341_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.815
cc_25 VNB N_VGND_c_384_n 0.0293274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_385_n 0.0280546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_386_n 0.0246411f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_28 VNB N_VGND_c_387_n 0.00749823f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.485
cc_29 VNB N_VGND_c_388_n 0.0189171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_389_n 0.0567269f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=2.055
cc_31 VNB N_VGND_c_390_n 0.275152f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=2.055
cc_32 VNB N_VGND_c_391_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.815
cc_33 VNB N_A_257_136#_c_423_n 0.00977457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_257_136#_c_424_n 0.00343423f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_35 VPB N_A_83_264#_c_70_n 0.0215842f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_36 VPB N_A_83_264#_c_65_n 0.00819876f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.542
cc_37 VPB N_A_83_264#_c_72_n 0.0103777f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.97
cc_38 VPB N_A_83_264#_c_73_n 0.00257348f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.815
cc_39 VPB N_A_83_264#_c_67_n 0.0028461f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=1.94
cc_40 VPB N_A_83_264#_c_75_n 0.0075506f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.14
cc_41 VPB N_A_83_264#_c_76_n 0.0346366f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.815
cc_42 VPB N_A_83_264#_c_77_n 0.00825296f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.105
cc_43 VPB N_A1_c_177_n 0.0192469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A1_c_175_n 0.0382181f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_45 VPB N_A1_c_176_n 0.00453552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A2_c_213_n 0.00741577f $X=-0.19 $Y=1.66 $X2=2.41 $Y2=1.96
cc_47 VPB N_A2_c_218_n 0.0215591f $X=-0.19 $Y=1.66 $X2=3.89 $Y2=1.96
cc_48 VPB N_B1_c_255_n 0.0180921f $X=-0.19 $Y=1.66 $X2=3.785 $Y2=0.68
cc_49 VPB B1 0.00109348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_B1_c_254_n 0.0322785f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_51 VPB N_C1_c_289_n 0.0489526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB C1 0.0090211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB X 0.0138434f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_54 VPB X 0.041687f $X=-0.19 $Y=1.66 $X2=2.395 $Y2=2.055
cc_55 VPB N_X_c_317_n 0.00779372f $X=-0.19 $Y=1.66 $X2=2.835 $Y2=1.235
cc_56 VPB N_VPWR_c_342_n 0.0149614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_343_n 0.03031f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.542
cc_58 VPB N_VPWR_c_344_n 0.0191515f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.14
cc_59 VPB N_VPWR_c_341_n 0.0668915f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.815
cc_60 VPB N_VPWR_c_346_n 0.0189171f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=1.235
cc_61 VPB N_VPWR_c_347_n 0.0398894f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.485
cc_62 VPB N_VPWR_c_348_n 0.0155543f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.485
cc_63 N_A_83_264#_c_66_n N_A1_M1002_g 7.84219e-19 $X=1.01 $Y=1.65 $X2=0 $Y2=0
cc_64 N_A_83_264#_c_68_n N_A1_M1002_g 0.00270451f $X=0.93 $Y=1.485 $X2=0 $Y2=0
cc_65 N_A_83_264#_c_80_p N_A1_c_177_n 0.0165434f $X=2.395 $Y=2.055 $X2=0 $Y2=0
cc_66 N_A_83_264#_c_73_n N_A1_c_177_n 0.00274859f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_67 N_A_83_264#_c_66_n N_A1_c_175_n 7.57698e-19 $X=1.01 $Y=1.65 $X2=0 $Y2=0
cc_68 N_A_83_264#_c_72_n N_A1_c_175_n 0.00369873f $X=1.01 $Y=1.97 $X2=0 $Y2=0
cc_69 N_A_83_264#_c_80_p N_A1_c_175_n 0.00334143f $X=2.395 $Y=2.055 $X2=0 $Y2=0
cc_70 N_A_83_264#_c_68_n N_A1_c_175_n 0.0101707f $X=0.93 $Y=1.485 $X2=0 $Y2=0
cc_71 N_A_83_264#_c_66_n N_A1_c_176_n 0.0114678f $X=1.01 $Y=1.65 $X2=0 $Y2=0
cc_72 N_A_83_264#_c_72_n N_A1_c_176_n 0.00916902f $X=1.01 $Y=1.97 $X2=0 $Y2=0
cc_73 N_A_83_264#_c_80_p N_A1_c_176_n 0.0466193f $X=2.395 $Y=2.055 $X2=0 $Y2=0
cc_74 N_A_83_264#_c_67_n N_A1_c_176_n 0.00919118f $X=2.75 $Y=1.94 $X2=0 $Y2=0
cc_75 N_A_83_264#_c_68_n N_A1_c_176_n 2.26109e-19 $X=0.93 $Y=1.485 $X2=0 $Y2=0
cc_76 N_A_83_264#_c_80_p N_A2_c_218_n 0.0137777f $X=2.395 $Y=2.055 $X2=0 $Y2=0
cc_77 N_A_83_264#_c_73_n N_A2_c_218_n 0.0146112f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_78 N_A_83_264#_c_67_n N_A2_c_218_n 0.00101779f $X=2.75 $Y=1.94 $X2=0 $Y2=0
cc_79 N_A_83_264#_c_77_n N_A2_c_218_n 0.00204153f $X=2.56 $Y=2.105 $X2=0 $Y2=0
cc_80 N_A_83_264#_c_67_n N_A2_M1006_g 0.00940242f $X=2.75 $Y=1.94 $X2=0 $Y2=0
cc_81 N_A_83_264#_c_96_p N_A2_M1006_g 0.00176342f $X=2.835 $Y=1.235 $X2=0 $Y2=0
cc_82 N_A_83_264#_c_97_p A2 0.0159143f $X=3.76 $Y=1.235 $X2=0 $Y2=0
cc_83 N_A_83_264#_c_73_n N_B1_c_255_n 0.0142372f $X=2.56 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_83_264#_c_67_n N_B1_c_255_n 0.00282452f $X=2.75 $Y=1.94 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_83_264#_c_100_p N_B1_c_255_n 0.00610156f $X=3.875 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_86 N_A_83_264#_c_77_n N_B1_c_255_n 0.00946578f $X=2.56 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_83_264#_c_67_n N_B1_M1004_g 0.00432432f $X=2.75 $Y=1.94 $X2=0 $Y2=0
cc_88 N_A_83_264#_c_97_p N_B1_M1004_g 0.0138851f $X=3.76 $Y=1.235 $X2=0 $Y2=0
cc_89 N_A_83_264#_c_69_n N_B1_M1004_g 0.00125475f $X=3.97 $Y=0.855 $X2=0 $Y2=0
cc_90 N_A_83_264#_c_67_n B1 0.0221103f $X=2.75 $Y=1.94 $X2=0 $Y2=0
cc_91 N_A_83_264#_c_97_p B1 0.0209068f $X=3.76 $Y=1.235 $X2=0 $Y2=0
cc_92 N_A_83_264#_c_100_p B1 0.0242484f $X=3.875 $Y=2.055 $X2=0 $Y2=0
cc_93 N_A_83_264#_c_67_n N_B1_c_254_n 0.0183725f $X=2.75 $Y=1.94 $X2=0 $Y2=0
cc_94 N_A_83_264#_c_97_p N_B1_c_254_n 0.00827816f $X=3.76 $Y=1.235 $X2=0 $Y2=0
cc_95 N_A_83_264#_c_100_p N_B1_c_254_n 0.0112314f $X=3.875 $Y=2.055 $X2=0 $Y2=0
cc_96 N_A_83_264#_c_97_p N_C1_M1000_g 0.00974156f $X=3.76 $Y=1.235 $X2=0 $Y2=0
cc_97 N_A_83_264#_c_69_n N_C1_M1000_g 0.0112161f $X=3.97 $Y=0.855 $X2=0 $Y2=0
cc_98 N_A_83_264#_c_100_p N_C1_c_289_n 0.0162082f $X=3.875 $Y=2.055 $X2=0 $Y2=0
cc_99 N_A_83_264#_c_75_n N_C1_c_289_n 0.00169682f $X=4.04 $Y=2.14 $X2=0 $Y2=0
cc_100 N_A_83_264#_c_76_n N_C1_c_289_n 0.014389f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_101 N_A_83_264#_c_69_n N_C1_c_289_n 0.00453775f $X=3.97 $Y=0.855 $X2=0 $Y2=0
cc_102 N_A_83_264#_c_97_p C1 0.00884799f $X=3.76 $Y=1.235 $X2=0 $Y2=0
cc_103 N_A_83_264#_c_100_p C1 0.015204f $X=3.875 $Y=2.055 $X2=0 $Y2=0
cc_104 N_A_83_264#_c_75_n C1 0.0246244f $X=4.04 $Y=2.14 $X2=0 $Y2=0
cc_105 N_A_83_264#_c_69_n C1 0.0286973f $X=3.97 $Y=0.855 $X2=0 $Y2=0
cc_106 N_A_83_264#_M1008_g N_X_c_315_n 0.00825483f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_83_264#_M1008_g N_X_c_316_n 0.00285209f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_83_264#_c_65_n N_X_c_316_n 2.24457e-19 $X=0.505 $Y=1.542 $X2=0 $Y2=0
cc_109 N_A_83_264#_c_124_p N_X_c_316_n 0.00138666f $X=0.93 $Y=1.485 $X2=0 $Y2=0
cc_110 N_A_83_264#_c_70_n X 0.00378032f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_83_264#_c_65_n X 6.90698e-19 $X=0.505 $Y=1.542 $X2=0 $Y2=0
cc_112 N_A_83_264#_c_72_n X 0.00516881f $X=1.01 $Y=1.97 $X2=0 $Y2=0
cc_113 N_A_83_264#_c_128_p X 0.00629613f $X=1.095 $Y=2.055 $X2=0 $Y2=0
cc_114 N_A_83_264#_c_124_p X 0.00153915f $X=0.93 $Y=1.485 $X2=0 $Y2=0
cc_115 N_A_83_264#_c_70_n X 0.0180242f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_83_264#_M1008_g N_X_c_317_n 0.00480212f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A_83_264#_c_65_n N_X_c_317_n 0.0116038f $X=0.505 $Y=1.542 $X2=0 $Y2=0
cc_118 N_A_83_264#_c_72_n N_X_c_317_n 0.00340852f $X=1.01 $Y=1.97 $X2=0 $Y2=0
cc_119 N_A_83_264#_c_124_p N_X_c_317_n 0.026181f $X=0.93 $Y=1.485 $X2=0 $Y2=0
cc_120 N_A_83_264#_c_72_n N_VPWR_M1005_d 5.52896e-19 $X=1.01 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_83_264#_c_80_p N_VPWR_M1005_d 0.0239925f $X=2.395 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_83_264#_c_128_p N_VPWR_M1005_d 0.00595103f $X=1.095 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_123 N_A_83_264#_c_100_p N_VPWR_M1003_d 0.0230282f $X=3.875 $Y=2.055 $X2=0
+ $Y2=0
cc_124 N_A_83_264#_c_73_n N_VPWR_c_342_n 0.0260221f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_125 N_A_83_264#_c_100_p N_VPWR_c_342_n 0.0623206f $X=3.875 $Y=2.055 $X2=0
+ $Y2=0
cc_126 N_A_83_264#_c_76_n N_VPWR_c_342_n 0.0260221f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_127 N_A_83_264#_c_73_n N_VPWR_c_343_n 0.014552f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_128 N_A_83_264#_c_76_n N_VPWR_c_344_n 0.0145938f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_129 N_A_83_264#_c_70_n N_VPWR_c_341_n 0.00865191f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_83_264#_c_73_n N_VPWR_c_341_n 0.0119791f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_131 N_A_83_264#_c_76_n N_VPWR_c_341_n 0.0120466f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_132 N_A_83_264#_c_70_n N_VPWR_c_346_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_83_264#_c_70_n N_VPWR_c_347_n 0.0183829f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A_83_264#_c_80_p N_VPWR_c_347_n 0.0567882f $X=2.395 $Y=2.055 $X2=0
+ $Y2=0
cc_135 N_A_83_264#_c_128_p N_VPWR_c_347_n 0.0151701f $X=1.095 $Y=2.055 $X2=0
+ $Y2=0
cc_136 N_A_83_264#_c_73_n N_VPWR_c_347_n 0.0206303f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_137 N_A_83_264#_c_124_p N_VPWR_c_347_n 0.00837395f $X=0.93 $Y=1.485 $X2=0
+ $Y2=0
cc_138 N_A_83_264#_c_68_n N_VPWR_c_347_n 0.00553603f $X=0.93 $Y=1.485 $X2=0
+ $Y2=0
cc_139 N_A_83_264#_c_80_p A_398_392# 0.00924457f $X=2.395 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_83_264#_M1008_g N_VGND_c_384_n 0.0198727f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_141 N_A_83_264#_c_66_n N_VGND_c_384_n 0.00155683f $X=1.01 $Y=1.65 $X2=0 $Y2=0
cc_142 N_A_83_264#_c_124_p N_VGND_c_384_n 0.0239345f $X=0.93 $Y=1.485 $X2=0
+ $Y2=0
cc_143 N_A_83_264#_c_68_n N_VGND_c_384_n 0.00727465f $X=0.93 $Y=1.485 $X2=0
+ $Y2=0
cc_144 N_A_83_264#_M1008_g N_VGND_c_388_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_83_264#_c_69_n N_VGND_c_389_n 0.00480029f $X=3.97 $Y=0.855 $X2=0
+ $Y2=0
cc_146 N_A_83_264#_M1008_g N_VGND_c_390_n 0.00828717f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_83_264#_c_69_n N_VGND_c_390_n 0.012096f $X=3.97 $Y=0.855 $X2=0 $Y2=0
cc_148 N_A_83_264#_c_97_p N_A_257_136#_M1006_d 0.00708637f $X=3.76 $Y=1.235
+ $X2=0 $Y2=0
cc_149 N_A_83_264#_c_96_p N_A_257_136#_M1006_d 0.00482969f $X=2.835 $Y=1.235
+ $X2=0 $Y2=0
cc_150 N_A_83_264#_c_80_p N_A_257_136#_c_427_n 0.00764285f $X=2.395 $Y=2.055
+ $X2=0 $Y2=0
cc_151 N_A_83_264#_c_96_p N_A_257_136#_c_427_n 0.0135241f $X=2.835 $Y=1.235
+ $X2=0 $Y2=0
cc_152 N_A_83_264#_c_77_n N_A_257_136#_c_427_n 0.00237837f $X=2.56 $Y=2.105
+ $X2=0 $Y2=0
cc_153 N_A_83_264#_M1008_g N_A_257_136#_c_424_n 0.00407387f $X=0.495 $Y=0.74
+ $X2=0 $Y2=0
cc_154 N_A_83_264#_c_80_p N_A_257_136#_c_424_n 0.00207755f $X=2.395 $Y=2.055
+ $X2=0 $Y2=0
cc_155 N_A_83_264#_c_97_p N_A_257_136#_c_432_n 0.02109f $X=3.76 $Y=1.235 $X2=0
+ $Y2=0
cc_156 N_A_83_264#_c_96_p N_A_257_136#_c_432_n 0.013831f $X=2.835 $Y=1.235 $X2=0
+ $Y2=0
cc_157 N_A_83_264#_c_69_n N_A_257_136#_c_432_n 0.00424382f $X=3.97 $Y=0.855
+ $X2=0 $Y2=0
cc_158 N_A_83_264#_c_97_p A_662_136# 0.00800139f $X=3.76 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A1_M1002_g N_A2_c_212_n 0.00187708f $X=1.69 $Y=1 $X2=-0.19 $Y2=-0.245
cc_160 N_A1_c_175_n N_A2_c_212_n 0.023699f $X=1.84 $Y=1.635 $X2=-0.19 $Y2=-0.245
cc_161 N_A1_c_176_n N_A2_c_212_n 0.00136073f $X=1.84 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A1_c_177_n N_A2_c_218_n 0.0538391f $X=1.915 $Y=1.885 $X2=0 $Y2=0
cc_163 N_A1_M1002_g N_A2_c_216_n 0.0129588f $X=1.69 $Y=1 $X2=0 $Y2=0
cc_164 N_A1_c_177_n N_VPWR_c_343_n 0.00413917f $X=1.915 $Y=1.885 $X2=0 $Y2=0
cc_165 N_A1_c_177_n N_VPWR_c_341_n 0.00812917f $X=1.915 $Y=1.885 $X2=0 $Y2=0
cc_166 N_A1_c_177_n N_VPWR_c_347_n 0.0177708f $X=1.915 $Y=1.885 $X2=0 $Y2=0
cc_167 N_A1_M1002_g N_VGND_c_384_n 0.00332473f $X=1.69 $Y=1 $X2=0 $Y2=0
cc_168 N_A1_M1002_g N_VGND_c_385_n 0.00385576f $X=1.69 $Y=1 $X2=0 $Y2=0
cc_169 N_A1_M1002_g N_VGND_c_386_n 0.00386669f $X=1.69 $Y=1 $X2=0 $Y2=0
cc_170 N_A1_M1002_g N_VGND_c_390_n 0.00454494f $X=1.69 $Y=1 $X2=0 $Y2=0
cc_171 N_A1_M1002_g N_A_257_136#_c_423_n 4.6447e-19 $X=1.69 $Y=1 $X2=0 $Y2=0
cc_172 N_A1_M1002_g N_A_257_136#_c_427_n 0.0136829f $X=1.69 $Y=1 $X2=0 $Y2=0
cc_173 N_A1_c_175_n N_A_257_136#_c_427_n 0.00154552f $X=1.84 $Y=1.635 $X2=0
+ $Y2=0
cc_174 N_A1_c_176_n N_A_257_136#_c_427_n 0.0271459f $X=1.84 $Y=1.635 $X2=0 $Y2=0
cc_175 N_A1_c_175_n N_A_257_136#_c_424_n 0.00191995f $X=1.84 $Y=1.635 $X2=0
+ $Y2=0
cc_176 N_A1_c_176_n N_A_257_136#_c_424_n 0.0197381f $X=1.84 $Y=1.635 $X2=0 $Y2=0
cc_177 N_A1_M1002_g N_A_257_136#_c_441_n 5.79196e-19 $X=1.69 $Y=1 $X2=0 $Y2=0
cc_178 N_A2_c_218_n N_B1_c_255_n 0.00843851f $X=2.335 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_179 A2 N_B1_M1004_g 0.0110521f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_180 N_A2_c_216_n N_B1_M1004_g 3.79406e-19 $X=2.49 $Y=0.405 $X2=0 $Y2=0
cc_181 N_A2_c_212_n N_B1_c_254_n 0.0182214f $X=2.335 $Y=1.5 $X2=0 $Y2=0
cc_182 A2 N_C1_M1000_g 0.00944212f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_183 N_A2_c_218_n N_VPWR_c_343_n 0.00445602f $X=2.335 $Y=1.885 $X2=0 $Y2=0
cc_184 N_A2_c_218_n N_VPWR_c_341_n 0.00858241f $X=2.335 $Y=1.885 $X2=0 $Y2=0
cc_185 N_A2_c_218_n N_VPWR_c_347_n 0.00246374f $X=2.335 $Y=1.885 $X2=0 $Y2=0
cc_186 A2 N_VGND_c_385_n 0.0325047f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_187 N_A2_c_216_n N_VGND_c_385_n 0.0147033f $X=2.49 $Y=0.405 $X2=0 $Y2=0
cc_188 A2 N_VGND_c_389_n 0.0938129f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_189 N_A2_c_216_n N_VGND_c_389_n 0.00730783f $X=2.49 $Y=0.405 $X2=0 $Y2=0
cc_190 A2 N_VGND_c_390_n 0.0517281f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_191 N_A2_c_216_n N_VGND_c_390_n 0.0105588f $X=2.49 $Y=0.405 $X2=0 $Y2=0
cc_192 N_A2_M1006_g N_A_257_136#_c_427_n 0.0145392f $X=2.35 $Y=1 $X2=0 $Y2=0
cc_193 N_A2_M1006_g N_A_257_136#_c_441_n 0.00443211f $X=2.35 $Y=1 $X2=0 $Y2=0
cc_194 N_A2_M1006_g N_A_257_136#_c_444_n 0.00477026f $X=2.35 $Y=1 $X2=0 $Y2=0
cc_195 A2 N_A_257_136#_c_444_n 0.0111303f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_196 N_A2_c_216_n N_A_257_136#_c_444_n 3.08235e-19 $X=2.49 $Y=0.405 $X2=0
+ $Y2=0
cc_197 A2 N_A_257_136#_c_432_n 0.050885f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_198 N_A2_c_216_n N_A_257_136#_c_432_n 9.34666e-19 $X=2.49 $Y=0.405 $X2=0
+ $Y2=0
cc_199 N_B1_M1004_g N_C1_M1000_g 0.0356518f $X=3.235 $Y=1 $X2=0 $Y2=0
cc_200 B1 N_C1_c_289_n 3.96013e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_201 N_B1_c_254_n N_C1_c_289_n 0.0140868f $X=3.17 $Y=1.635 $X2=0 $Y2=0
cc_202 B1 C1 0.0153874f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_203 N_B1_c_254_n C1 3.90152e-19 $X=3.17 $Y=1.635 $X2=0 $Y2=0
cc_204 N_B1_c_255_n N_VPWR_c_342_n 0.0183824f $X=2.785 $Y=1.885 $X2=0 $Y2=0
cc_205 N_B1_c_255_n N_VPWR_c_343_n 0.00445602f $X=2.785 $Y=1.885 $X2=0 $Y2=0
cc_206 N_B1_c_255_n N_VPWR_c_341_n 0.00861803f $X=2.785 $Y=1.885 $X2=0 $Y2=0
cc_207 N_B1_M1004_g N_VGND_c_389_n 4.78105e-19 $X=3.235 $Y=1 $X2=0 $Y2=0
cc_208 N_B1_M1004_g N_A_257_136#_c_427_n 9.56449e-19 $X=3.235 $Y=1 $X2=0 $Y2=0
cc_209 N_B1_M1004_g N_A_257_136#_c_441_n 0.00194622f $X=3.235 $Y=1 $X2=0 $Y2=0
cc_210 N_B1_M1004_g N_A_257_136#_c_432_n 0.00380359f $X=3.235 $Y=1 $X2=0 $Y2=0
cc_211 N_B1_c_254_n N_A_257_136#_c_432_n 8.28061e-19 $X=3.17 $Y=1.635 $X2=0
+ $Y2=0
cc_212 N_C1_c_289_n N_VPWR_c_342_n 0.0183824f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_213 N_C1_c_289_n N_VPWR_c_344_n 0.00445602f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_214 N_C1_c_289_n N_VPWR_c_341_n 0.00865213f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_215 N_C1_M1000_g N_VGND_c_389_n 0.00206323f $X=3.71 $Y=1 $X2=0 $Y2=0
cc_216 N_C1_M1000_g N_VGND_c_390_n 0.00212097f $X=3.71 $Y=1 $X2=0 $Y2=0
cc_217 N_C1_M1000_g N_A_257_136#_c_432_n 5.49226e-19 $X=3.71 $Y=1 $X2=0 $Y2=0
cc_218 X N_VPWR_c_341_n 0.0131546f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_219 X N_VPWR_c_346_n 0.0159324f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_220 X N_VPWR_c_347_n 0.0264456f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_221 N_X_c_315_n N_VGND_c_384_n 0.0312028f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_222 N_X_c_315_n N_VGND_c_388_n 0.0159025f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_223 N_X_c_315_n N_VGND_c_390_n 0.0131064f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_224 N_VGND_c_384_n N_A_257_136#_c_423_n 0.0252292f $X=0.78 $Y=0.515 $X2=0
+ $Y2=0
cc_225 N_VGND_c_385_n N_A_257_136#_c_423_n 0.0120549f $X=1.96 $Y=0.84 $X2=0
+ $Y2=0
cc_226 N_VGND_c_386_n N_A_257_136#_c_423_n 0.00628283f $X=1.765 $Y=0 $X2=0 $Y2=0
cc_227 N_VGND_c_390_n N_A_257_136#_c_423_n 0.00974349f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_M1002_d N_A_257_136#_c_427_n 0.0136241f $X=1.765 $Y=0.68 $X2=0
+ $Y2=0
cc_229 N_VGND_c_385_n N_A_257_136#_c_427_n 0.0234958f $X=1.96 $Y=0.84 $X2=0
+ $Y2=0
cc_230 N_VGND_c_385_n N_A_257_136#_c_444_n 0.00959329f $X=1.96 $Y=0.84 $X2=0
+ $Y2=0
