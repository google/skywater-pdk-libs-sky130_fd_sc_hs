* File: sky130_fd_sc_hs__ebufn_8.pex.spice
* Created: Thu Aug 27 20:44:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__EBUFN_8%A_84_48# 1 2 9 11 13 16 18 20 23 25 27 30 32
+ 34 37 39 41 44 46 48 49 51 54 56 58 61 63 68 71 72 73 74 79 82 84 86 88 90 91
+ 93 98 102 120
c272 97 0 6.69633e-20 $X=3.655 $Y=1.485
c273 71 0 8.42804e-20 $X=3.955 $Y=2.05
c274 61 0 1.9142e-19 $X=3.81 $Y=0.74
c275 56 0 1.85036e-19 $X=3.795 $Y=1.765
r276 120 121 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=3.795 $Y=1.542
+ $X2=3.81 $Y2=1.542
r277 117 118 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=3.31 $Y=1.542
+ $X2=3.325 $Y2=1.542
r278 116 117 63.9257 $w=3.77e-07 $l=5e-07 $layer=POLY_cond $X=2.81 $Y=1.542
+ $X2=3.31 $Y2=1.542
r279 115 116 57.5332 $w=3.77e-07 $l=4.5e-07 $layer=POLY_cond $X=2.36 $Y=1.542
+ $X2=2.81 $Y2=1.542
r280 114 115 6.39257 $w=3.77e-07 $l=5e-08 $layer=POLY_cond $X=2.31 $Y=1.542
+ $X2=2.36 $Y2=1.542
r281 113 114 51.1406 $w=3.77e-07 $l=4e-07 $layer=POLY_cond $X=1.91 $Y=1.542
+ $X2=2.31 $Y2=1.542
r282 112 113 12.7851 $w=3.77e-07 $l=1e-07 $layer=POLY_cond $X=1.81 $Y=1.542
+ $X2=1.91 $Y2=1.542
r283 111 112 51.1406 $w=3.77e-07 $l=4e-07 $layer=POLY_cond $X=1.41 $Y=1.542
+ $X2=1.81 $Y2=1.542
r284 110 111 3.83554 $w=3.77e-07 $l=3e-08 $layer=POLY_cond $X=1.38 $Y=1.542
+ $X2=1.41 $Y2=1.542
r285 107 108 4.4748 $w=3.77e-07 $l=3.5e-08 $layer=POLY_cond $X=0.925 $Y=1.542
+ $X2=0.96 $Y2=1.542
r286 106 107 53.0584 $w=3.77e-07 $l=4.15e-07 $layer=POLY_cond $X=0.51 $Y=1.542
+ $X2=0.925 $Y2=1.542
r287 105 106 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.542
+ $X2=0.51 $Y2=1.542
r288 98 100 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.67 $Y=2.135
+ $X2=7.67 $Y2=2.305
r289 96 120 35.1592 $w=3.77e-07 $l=2.75e-07 $layer=POLY_cond $X=3.52 $Y=1.542
+ $X2=3.795 $Y2=1.542
r290 96 118 24.931 $w=3.77e-07 $l=1.95e-07 $layer=POLY_cond $X=3.52 $Y=1.542
+ $X2=3.325 $Y2=1.542
r291 95 97 7.4145 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.52 $Y=1.485
+ $X2=3.655 $Y2=1.485
r292 95 96 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=3.52
+ $Y=1.485 $X2=3.52 $Y2=1.485
r293 92 93 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=10.23 $Y=1.01
+ $X2=10.23 $Y2=1.72
r294 90 93 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.145 $Y=1.805
+ $X2=10.23 $Y2=1.72
r295 90 91 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=10.145 $Y=1.805
+ $X2=9.945 $Y2=1.805
r296 89 104 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.93 $Y=0.925
+ $X2=9.805 $Y2=0.925
r297 88 92 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.145 $Y=0.925
+ $X2=10.23 $Y2=1.01
r298 88 89 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.145 $Y=0.925
+ $X2=9.93 $Y2=0.925
r299 84 104 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.805 $Y=0.84
+ $X2=9.805 $Y2=0.925
r300 84 86 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=9.805 $Y=0.84
+ $X2=9.805 $Y2=0.505
r301 80 102 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.805 $Y=2.39
+ $X2=9.805 $Y2=2.305
r302 80 82 17.4924 $w=2.78e-07 $l=4.25e-07 $layer=LI1_cond $X=9.805 $Y=2.39
+ $X2=9.805 $Y2=2.815
r303 77 102 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.805 $Y=2.22
+ $X2=9.805 $Y2=2.305
r304 77 79 9.67229 $w=2.78e-07 $l=2.35e-07 $layer=LI1_cond $X=9.805 $Y=2.22
+ $X2=9.805 $Y2=1.985
r305 76 91 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=9.805 $Y=1.89
+ $X2=9.945 $Y2=1.805
r306 76 79 3.91007 $w=2.78e-07 $l=9.5e-08 $layer=LI1_cond $X=9.805 $Y=1.89
+ $X2=9.805 $Y2=1.985
r307 75 100 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=2.305
+ $X2=7.67 $Y2=2.305
r308 74 102 3.18746 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=9.665 $Y=2.305
+ $X2=9.805 $Y2=2.305
r309 74 75 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=9.665 $Y=2.305
+ $X2=7.755 $Y2=2.305
r310 72 98 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=2.135
+ $X2=7.67 $Y2=2.135
r311 72 73 231.278 $w=1.68e-07 $l=3.545e-06 $layer=LI1_cond $X=7.585 $Y=2.135
+ $X2=4.04 $Y2=2.135
r312 71 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.955 $Y=2.05
+ $X2=4.04 $Y2=2.135
r313 70 71 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.955 $Y=1.65
+ $X2=3.955 $Y2=2.05
r314 68 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.87 $Y=1.565
+ $X2=3.955 $Y2=1.65
r315 68 97 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.87 $Y=1.565
+ $X2=3.655 $Y2=1.565
r316 66 110 30.6844 $w=3.77e-07 $l=2.4e-07 $layer=POLY_cond $X=1.14 $Y=1.542
+ $X2=1.38 $Y2=1.542
r317 66 108 23.0133 $w=3.77e-07 $l=1.8e-07 $layer=POLY_cond $X=1.14 $Y=1.542
+ $X2=0.96 $Y2=1.542
r318 65 66 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=1.14
+ $Y=1.485 $X2=1.14 $Y2=1.485
r319 63 95 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=3.49 $Y=1.485
+ $X2=3.52 $Y2=1.485
r320 63 65 82.0679 $w=3.28e-07 $l=2.35e-06 $layer=LI1_cond $X=3.49 $Y=1.485
+ $X2=1.14 $Y2=1.485
r321 59 121 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.81 $Y=1.32
+ $X2=3.81 $Y2=1.542
r322 59 61 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.81 $Y=1.32
+ $X2=3.81 $Y2=0.74
r323 56 120 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.795 $Y=1.765
+ $X2=3.795 $Y2=1.542
r324 56 58 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.795 $Y=1.765
+ $X2=3.795 $Y2=2.4
r325 52 118 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.325 $Y=1.32
+ $X2=3.325 $Y2=1.542
r326 52 54 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.325 $Y=1.32
+ $X2=3.325 $Y2=0.74
r327 49 117 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.31 $Y=1.765
+ $X2=3.31 $Y2=1.542
r328 49 51 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.31 $Y=1.765
+ $X2=3.31 $Y2=2.4
r329 46 116 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.81 $Y=1.765
+ $X2=2.81 $Y2=1.542
r330 46 48 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.81 $Y=1.765
+ $X2=2.81 $Y2=2.4
r331 42 116 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.81 $Y=1.32
+ $X2=2.81 $Y2=1.542
r332 42 44 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.81 $Y=1.32
+ $X2=2.81 $Y2=0.74
r333 39 115 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=1.542
r334 39 41 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=2.4
r335 35 114 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.31 $Y=1.32
+ $X2=2.31 $Y2=1.542
r336 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.31 $Y=1.32
+ $X2=2.31 $Y2=0.74
r337 32 113 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=1.542
r338 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=2.4
r339 28 112 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.81 $Y=1.32
+ $X2=1.81 $Y2=1.542
r340 28 30 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.81 $Y=1.32
+ $X2=1.81 $Y2=0.74
r341 25 111 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=1.542
r342 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=2.4
r343 21 110 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.38 $Y=1.32
+ $X2=1.38 $Y2=1.542
r344 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.38 $Y=1.32
+ $X2=1.38 $Y2=0.74
r345 18 108 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.542
r346 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r347 14 107 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.925 $Y=1.32
+ $X2=0.925 $Y2=1.542
r348 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.925 $Y=1.32
+ $X2=0.925 $Y2=0.74
r349 11 106 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.542
r350 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r351 7 105 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=1.542
r352 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.74
r353 2 82 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.84 $X2=9.83 $Y2=2.815
r354 2 79 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.84 $X2=9.83 $Y2=1.985
r355 1 104 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=9.705
+ $Y=0.37 $X2=9.845 $Y2=0.925
r356 1 86 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=9.705
+ $Y=0.37 $X2=9.845 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_8%A_833_48# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 24 25 27 29 30 32 34 35 37 39 40 42 44 45 48 49 50 51 52 53 54 55 56 58 59 62
+ 64 66 68
c165 58 0 1.51364e-19 $X=8.01 $Y=1.8
c166 17 0 2.61838e-20 $X=5.1 $Y=1.185
c167 11 0 6.69633e-20 $X=4.315 $Y=1.26
c168 7 0 7.54658e-20 $X=4.24 $Y=1.185
r169 71 73 3.15083 $w=4.84e-07 $l=1.25e-07 $layer=LI1_cond $X=7.885 $Y=0.67
+ $X2=8.01 $Y2=0.67
r170 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.885
+ $Y=0.505 $X2=7.885 $Y2=0.505
r171 66 68 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=8.095 $Y=1.925
+ $X2=8.77 $Y2=1.925
r172 62 72 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=8.565 $Y=0.505
+ $X2=7.885 $Y2=0.505
r173 61 64 7.49781 $w=6.68e-07 $l=4.2e-07 $layer=LI1_cond $X=8.565 $Y=0.675
+ $X2=8.985 $Y2=0.675
r174 61 62 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.565
+ $Y=0.505 $X2=8.565 $Y2=0.505
r175 59 73 2.5084 $w=6.7e-07 $l=8.74643e-08 $layer=LI1_cond $X=8.095 $Y=0.675
+ $X2=8.01 $Y2=0.67
r176 59 61 8.3904 $w=6.68e-07 $l=4.7e-07 $layer=LI1_cond $X=8.095 $Y=0.675
+ $X2=8.565 $Y2=0.675
r177 58 66 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.01 $Y=1.8
+ $X2=8.095 $Y2=1.925
r178 57 73 6.95298 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=8.01 $Y=1.01
+ $X2=8.01 $Y2=0.67
r179 57 58 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.01 $Y=1.01
+ $X2=8.01 $Y2=1.8
r180 56 72 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.87 $Y=0.505
+ $X2=7.885 $Y2=0.505
r181 47 56 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.795 $Y=0.67
+ $X2=7.87 $Y2=0.505
r182 47 48 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=7.795 $Y=0.67
+ $X2=7.795 $Y2=1.185
r183 46 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.325 $Y=1.26
+ $X2=7.25 $Y2=1.26
r184 45 48 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.72 $Y=1.26
+ $X2=7.795 $Y2=1.185
r185 45 46 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.72 $Y=1.26
+ $X2=7.325 $Y2=1.26
r186 42 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.25 $Y=1.185
+ $X2=7.25 $Y2=1.26
r187 42 44 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.25 $Y=1.185
+ $X2=7.25 $Y2=0.74
r188 41 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.895 $Y=1.26
+ $X2=6.82 $Y2=1.26
r189 40 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.175 $Y=1.26
+ $X2=7.25 $Y2=1.26
r190 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.175 $Y=1.26
+ $X2=6.895 $Y2=1.26
r191 37 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.82 $Y=1.185
+ $X2=6.82 $Y2=1.26
r192 37 39 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.82 $Y=1.185
+ $X2=6.82 $Y2=0.74
r193 36 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.465 $Y=1.26
+ $X2=6.39 $Y2=1.26
r194 35 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.745 $Y=1.26
+ $X2=6.82 $Y2=1.26
r195 35 36 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.745 $Y=1.26
+ $X2=6.465 $Y2=1.26
r196 32 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.39 $Y=1.185
+ $X2=6.39 $Y2=1.26
r197 32 34 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.39 $Y=1.185
+ $X2=6.39 $Y2=0.74
r198 31 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.035 $Y=1.26
+ $X2=5.96 $Y2=1.26
r199 30 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.315 $Y=1.26
+ $X2=6.39 $Y2=1.26
r200 30 31 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.315 $Y=1.26
+ $X2=6.035 $Y2=1.26
r201 27 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.96 $Y=1.185
+ $X2=5.96 $Y2=1.26
r202 27 29 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.96 $Y=1.185
+ $X2=5.96 $Y2=0.74
r203 26 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.605 $Y=1.26
+ $X2=5.53 $Y2=1.26
r204 25 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.885 $Y=1.26
+ $X2=5.96 $Y2=1.26
r205 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.885 $Y=1.26
+ $X2=5.605 $Y2=1.26
r206 22 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.53 $Y=1.185
+ $X2=5.53 $Y2=1.26
r207 22 24 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.53 $Y=1.185
+ $X2=5.53 $Y2=0.74
r208 21 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.175 $Y=1.26
+ $X2=5.1 $Y2=1.26
r209 20 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.455 $Y=1.26
+ $X2=5.53 $Y2=1.26
r210 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.455 $Y=1.26
+ $X2=5.175 $Y2=1.26
r211 17 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.1 $Y=1.185
+ $X2=5.1 $Y2=1.26
r212 17 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.1 $Y=1.185
+ $X2=5.1 $Y2=0.74
r213 16 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.745 $Y=1.26
+ $X2=4.67 $Y2=1.26
r214 15 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.025 $Y=1.26
+ $X2=5.1 $Y2=1.26
r215 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.025 $Y=1.26
+ $X2=4.745 $Y2=1.26
r216 12 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.67 $Y=1.185
+ $X2=4.67 $Y2=1.26
r217 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.67 $Y=1.185
+ $X2=4.67 $Y2=0.74
r218 10 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.595 $Y=1.26
+ $X2=4.67 $Y2=1.26
r219 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.595 $Y=1.26
+ $X2=4.315 $Y2=1.26
r220 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.24 $Y=1.185
+ $X2=4.315 $Y2=1.26
r221 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.24 $Y=1.185
+ $X2=4.24 $Y2=0.74
r222 2 68 600 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=8.52
+ $Y=1.84 $X2=8.77 $Y2=1.965
r223 1 64 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=8.84
+ $Y=0.37 $X2=8.985 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_8%TE_B 1 3 4 5 6 8 9 11 13 14 16 18 19 21 23
+ 24 26 28 29 31 33 34 36 38 41 42 43 45 46 48 49 50 51 52 53 54 55 56 57 58 65
+ 67
c184 31 0 1.51364e-19 $X=7.26 $Y=1.765
r185 67 68 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.11
+ $Y=1.385 $X2=9.11 $Y2=1.385
r186 63 65 47.8511 $w=5.45e-07 $l=1.65e-07 $layer=POLY_cond $X=8.43 $Y=1.492
+ $X2=8.265 $Y2=1.492
r187 63 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.43
+ $Y=1.385 $X2=8.43 $Y2=1.385
r188 58 68 7.78678 $w=3.68e-07 $l=2.5e-07 $layer=LI1_cond $X=9.36 $Y=1.365
+ $X2=9.11 $Y2=1.365
r189 57 68 7.16384 $w=3.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=9.11 $Y2=1.365
r190 57 64 14.0162 $w=3.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=8.43 $Y2=1.365
r191 56 64 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=8.4 $Y=1.365
+ $X2=8.43 $Y2=1.365
r192 46 67 50.4302 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.2 $Y=1.22
+ $X2=9.03 $Y2=1.22
r193 46 48 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.2 $Y=1.22 $X2=9.2
+ $Y2=0.74
r194 43 67 50.4302 $w=1.5e-07 $l=5.81292e-07 $layer=POLY_cond $X=9.105 $Y=1.765
+ $X2=9.03 $Y2=1.22
r195 43 45 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.105 $Y=1.765
+ $X2=9.105 $Y2=2.4
r196 42 63 10.5042 $w=5.45e-07 $l=1.07e-07 $layer=POLY_cond $X=8.537 $Y=1.492
+ $X2=8.43 $Y2=1.492
r197 41 67 10.2225 $w=5.45e-07 $l=2.72e-07 $layer=POLY_cond $X=9.03 $Y=1.492
+ $X2=9.03 $Y2=1.22
r198 41 42 48.3981 $w=5.45e-07 $l=4.93e-07 $layer=POLY_cond $X=9.03 $Y=1.492
+ $X2=8.537 $Y2=1.492
r199 40 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.955 $Y=1.69
+ $X2=7.88 $Y2=1.69
r200 40 65 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.955 $Y=1.69
+ $X2=8.265 $Y2=1.69
r201 36 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.88 $Y=1.765
+ $X2=7.88 $Y2=1.69
r202 36 38 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.88 $Y=1.765
+ $X2=7.88 $Y2=2.4
r203 35 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.335 $Y=1.69
+ $X2=7.26 $Y2=1.69
r204 34 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.805 $Y=1.69
+ $X2=7.88 $Y2=1.69
r205 34 35 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=7.805 $Y=1.69 $X2=7.335
+ $Y2=1.69
r206 31 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.26 $Y=1.765
+ $X2=7.26 $Y2=1.69
r207 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.26 $Y=1.765
+ $X2=7.26 $Y2=2.4
r208 30 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.885 $Y=1.69
+ $X2=6.81 $Y2=1.69
r209 29 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.185 $Y=1.69
+ $X2=7.26 $Y2=1.69
r210 29 30 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=7.185 $Y=1.69
+ $X2=6.885 $Y2=1.69
r211 26 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.81 $Y=1.765
+ $X2=6.81 $Y2=1.69
r212 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.81 $Y=1.765
+ $X2=6.81 $Y2=2.4
r213 25 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.335 $Y=1.69
+ $X2=6.26 $Y2=1.69
r214 24 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.735 $Y=1.69
+ $X2=6.81 $Y2=1.69
r215 24 25 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.735 $Y=1.69
+ $X2=6.335 $Y2=1.69
r216 21 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.26 $Y=1.765
+ $X2=6.26 $Y2=1.69
r217 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.26 $Y=1.765
+ $X2=6.26 $Y2=2.4
r218 20 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.885 $Y=1.69
+ $X2=5.81 $Y2=1.69
r219 19 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.185 $Y=1.69
+ $X2=6.26 $Y2=1.69
r220 19 20 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=6.185 $Y=1.69
+ $X2=5.885 $Y2=1.69
r221 16 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.81 $Y=1.765
+ $X2=5.81 $Y2=1.69
r222 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.81 $Y=1.765
+ $X2=5.81 $Y2=2.4
r223 15 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.335 $Y=1.69
+ $X2=5.26 $Y2=1.69
r224 14 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.735 $Y=1.69
+ $X2=5.81 $Y2=1.69
r225 14 15 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.735 $Y=1.69
+ $X2=5.335 $Y2=1.69
r226 11 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.26 $Y=1.765
+ $X2=5.26 $Y2=1.69
r227 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.26 $Y=1.765
+ $X2=5.26 $Y2=2.4
r228 10 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.885 $Y=1.69
+ $X2=4.81 $Y2=1.69
r229 9 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.185 $Y=1.69
+ $X2=5.26 $Y2=1.69
r230 9 10 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=5.185 $Y=1.69 $X2=4.885
+ $Y2=1.69
r231 6 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.81 $Y=1.765
+ $X2=4.81 $Y2=1.69
r232 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.81 $Y=1.765
+ $X2=4.81 $Y2=2.4
r233 4 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.735 $Y=1.69
+ $X2=4.81 $Y2=1.69
r234 4 5 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.735 $Y=1.69 $X2=4.335
+ $Y2=1.69
r235 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.26 $Y=1.765
+ $X2=4.335 $Y2=1.69
r236 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.26 $Y=1.765
+ $X2=4.26 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_8%A 1 3 4 6 7 9 10 12 13 20
r50 20 21 0.533186 $w=4.52e-07 $l=5e-09 $layer=POLY_cond $X=10.055 $Y=1.492
+ $X2=10.06 $Y2=1.492
r51 18 20 26.1261 $w=4.52e-07 $l=2.45e-07 $layer=POLY_cond $X=9.81 $Y=1.492
+ $X2=10.055 $Y2=1.492
r52 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.81
+ $Y=1.385 $X2=9.81 $Y2=1.385
r53 16 18 19.1947 $w=4.52e-07 $l=1.8e-07 $layer=POLY_cond $X=9.63 $Y=1.492
+ $X2=9.81 $Y2=1.492
r54 15 16 2.66593 $w=4.52e-07 $l=2.5e-08 $layer=POLY_cond $X=9.605 $Y=1.492
+ $X2=9.63 $Y2=1.492
r55 13 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.81 $Y=1.295 $X2=9.81
+ $Y2=1.385
r56 10 21 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=10.06 $Y=1.22
+ $X2=10.06 $Y2=1.492
r57 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.06 $Y=1.22
+ $X2=10.06 $Y2=0.74
r58 7 20 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=10.055 $Y=1.765
+ $X2=10.055 $Y2=1.492
r59 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.055 $Y=1.765
+ $X2=10.055 $Y2=2.4
r60 4 16 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=9.63 $Y=1.22 $X2=9.63
+ $Y2=1.492
r61 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.63 $Y=1.22 $X2=9.63
+ $Y2=0.74
r62 1 15 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=9.605 $Y=1.765
+ $X2=9.605 $Y2=1.492
r63 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.605 $Y=1.765
+ $X2=9.605 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_8%A_28_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 40
+ 44 46 50 52 54 55 56 60 64 66 68 69 70 74 76 79 82
r138 82 85 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=8.105 $Y=2.645
+ $X2=8.105 $Y2=2.77
r139 79 80 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.035 $Y=2.475
+ $X2=7.035 $Y2=2.645
r140 67 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.2 $Y=2.645
+ $X2=7.035 $Y2=2.645
r141 66 82 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.94 $Y=2.645
+ $X2=8.105 $Y2=2.645
r142 66 67 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=7.94 $Y=2.645
+ $X2=7.2 $Y2=2.645
r143 65 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.2 $Y=2.475
+ $X2=6.035 $Y2=2.475
r144 64 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=2.475
+ $X2=7.035 $Y2=2.475
r145 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.87 $Y=2.475
+ $X2=6.2 $Y2=2.475
r146 61 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.2 $Y=2.475
+ $X2=5.035 $Y2=2.475
r147 60 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.87 $Y=2.475
+ $X2=6.035 $Y2=2.475
r148 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.87 $Y=2.475
+ $X2=5.2 $Y2=2.475
r149 57 72 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=2.475
+ $X2=4.035 $Y2=2.475
r150 56 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.87 $Y=2.475
+ $X2=5.035 $Y2=2.475
r151 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.87 $Y=2.475
+ $X2=4.2 $Y2=2.475
r152 54 72 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=2.56
+ $X2=4.035 $Y2=2.475
r153 54 55 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.035 $Y=2.56
+ $X2=4.035 $Y2=2.905
r154 53 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.19 $Y=2.99
+ $X2=3.055 $Y2=2.99
r155 52 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.87 $Y=2.99
+ $X2=4.035 $Y2=2.905
r156 52 53 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.87 $Y=2.99
+ $X2=3.19 $Y2=2.99
r157 48 70 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=2.905
+ $X2=3.055 $Y2=2.99
r158 48 50 24.7562 $w=2.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.055 $Y=2.905
+ $X2=3.055 $Y2=2.325
r159 47 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=2.99
+ $X2=2.135 $Y2=2.99
r160 46 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.92 $Y=2.99
+ $X2=3.055 $Y2=2.99
r161 46 47 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.92 $Y=2.99 $X2=2.22
+ $Y2=2.99
r162 42 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=2.905
+ $X2=2.135 $Y2=2.99
r163 42 44 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.135 $Y=2.905
+ $X2=2.135 $Y2=2.325
r164 41 68 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.35 $Y=2.99
+ $X2=1.217 $Y2=2.99
r165 40 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=2.99
+ $X2=2.135 $Y2=2.99
r166 40 41 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.05 $Y=2.99 $X2=1.35
+ $Y2=2.99
r167 36 68 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.217 $Y=2.905
+ $X2=1.217 $Y2=2.99
r168 36 38 25.2233 $w=2.63e-07 $l=5.8e-07 $layer=LI1_cond $X=1.217 $Y=2.905
+ $X2=1.217 $Y2=2.325
r169 34 68 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.217 $Y2=2.99
r170 34 35 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.37 $Y2=2.99
r171 30 33 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.245 $Y=1.985
+ $X2=0.245 $Y2=2.815
r172 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.245 $Y=2.905
+ $X2=0.37 $Y2=2.99
r173 28 33 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.245 $Y=2.905
+ $X2=0.245 $Y2=2.815
r174 9 85 600 $w=1.7e-07 $l=1.0022e-06 $layer=licon1_PDIFF $count=1 $X=7.955
+ $Y=1.84 $X2=8.105 $Y2=2.77
r175 8 79 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=6.885
+ $Y=1.84 $X2=7.035 $Y2=2.475
r176 7 76 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=5.885
+ $Y=1.84 $X2=6.035 $Y2=2.475
r177 6 74 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=4.885
+ $Y=1.84 $X2=5.035 $Y2=2.475
r178 5 72 300 $w=1.7e-07 $l=7.12741e-07 $layer=licon1_PDIFF $count=2 $X=3.87
+ $Y=1.84 $X2=4.035 $Y2=2.475
r179 4 50 300 $w=1.7e-07 $l=5.7639e-07 $layer=licon1_PDIFF $count=2 $X=2.885
+ $Y=1.84 $X2=3.085 $Y2=2.325
r180 3 44 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=1.985
+ $Y=1.84 $X2=2.135 $Y2=2.325
r181 2 38 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.325
r182 1 33 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r183 1 30 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_8%Z 1 2 3 4 5 6 7 8 27 29 31 35 39 41 43 47 51
+ 53 55 57 59 63 67 68 70 72 73 76 77 78 85 89
c133 57 0 1.85036e-19 $X=3.535 $Y=1.99
c134 55 0 5.58653e-20 $X=3.43 $Y=1.065
r135 83 89 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.71 $Y=0.98
+ $X2=0.71 $Y2=0.925
r136 77 78 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=1.295
+ $X2=0.69 $Y2=1.665
r137 77 90 5.76222 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=0.69 $Y=1.295
+ $X2=0.69 $Y2=1.15
r138 76 83 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.065
+ $X2=0.71 $Y2=0.98
r139 76 90 3.05675 $w=3.1e-07 $l=9.44722e-08 $layer=LI1_cond $X=0.71 $Y=1.065
+ $X2=0.69 $Y2=1.15
r140 76 89 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.71 $Y=0.91
+ $X2=0.71 $Y2=0.925
r141 76 85 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.71 $Y=0.91
+ $X2=0.71 $Y2=0.76
r142 65 78 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=0.69 $Y=1.82
+ $X2=0.69 $Y2=1.665
r143 65 67 2.94878 $w=3.22e-07 $l=9.97246e-08 $layer=LI1_cond $X=0.69 $Y=1.82
+ $X2=0.722 $Y2=1.905
r144 61 63 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.595 $Y=0.98
+ $X2=3.595 $Y2=0.76
r145 57 75 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=1.99
+ $X2=3.535 $Y2=1.905
r146 57 59 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=3.535 $Y=1.99
+ $X2=3.535 $Y2=2.65
r147 56 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=1.065
+ $X2=2.595 $Y2=1.065
r148 55 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.43 $Y=1.065
+ $X2=3.595 $Y2=0.98
r149 55 56 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.43 $Y=1.065
+ $X2=2.76 $Y2=1.065
r150 54 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=1.905
+ $X2=2.585 $Y2=1.905
r151 53 75 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.37 $Y=1.905
+ $X2=3.535 $Y2=1.905
r152 53 54 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.37 $Y=1.905
+ $X2=2.75 $Y2=1.905
r153 49 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.98
+ $X2=2.595 $Y2=1.065
r154 49 51 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.595 $Y=0.98
+ $X2=2.595 $Y2=0.76
r155 45 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=1.99
+ $X2=2.585 $Y2=1.905
r156 45 47 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=2.585 $Y=1.99
+ $X2=2.585 $Y2=2.65
r157 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=1.905
+ $X2=1.685 $Y2=1.905
r158 43 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=1.905
+ $X2=2.585 $Y2=1.905
r159 43 44 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.42 $Y=1.905
+ $X2=1.85 $Y2=1.905
r160 42 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.76 $Y=1.065
+ $X2=1.595 $Y2=1.065
r161 41 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=1.065
+ $X2=2.595 $Y2=1.065
r162 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.43 $Y=1.065
+ $X2=1.76 $Y2=1.065
r163 37 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=1.99
+ $X2=1.685 $Y2=1.905
r164 37 39 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=1.685 $Y=1.99
+ $X2=1.685 $Y2=2.65
r165 33 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.595 $Y=0.98
+ $X2=1.595 $Y2=1.065
r166 33 35 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.595 $Y=0.98
+ $X2=1.595 $Y2=0.76
r167 32 67 3.72223 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.9 $Y=1.905
+ $X2=0.722 $Y2=1.905
r168 31 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=1.905
+ $X2=1.685 $Y2=1.905
r169 31 32 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.52 $Y=1.905
+ $X2=0.9 $Y2=1.905
r170 30 76 3.57226 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=1.065
+ $X2=0.71 $Y2=1.065
r171 29 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.43 $Y=1.065
+ $X2=1.595 $Y2=1.065
r172 29 30 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.43 $Y=1.065
+ $X2=0.875 $Y2=1.065
r173 25 67 2.94878 $w=3.22e-07 $l=8.5e-08 $layer=LI1_cond $X=0.722 $Y=1.99
+ $X2=0.722 $Y2=1.905
r174 25 27 21.4257 $w=3.53e-07 $l=6.6e-07 $layer=LI1_cond $X=0.722 $Y=1.99
+ $X2=0.722 $Y2=2.65
r175 8 75 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.84 $X2=3.535 $Y2=1.97
r176 8 59 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.84 $X2=3.535 $Y2=2.65
r177 7 72 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.84 $X2=2.585 $Y2=1.97
r178 7 47 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.84 $X2=2.585 $Y2=2.65
r179 6 70 400 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.685 $Y2=1.97
r180 6 39 400 $w=1.7e-07 $l=9.04489e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.685 $Y2=2.65
r181 5 67 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=1.97
r182 5 27 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.65
r183 4 63 182 $w=1.7e-07 $l=4.77651e-07 $layer=licon1_NDIFF $count=1 $X=3.4
+ $Y=0.37 $X2=3.595 $Y2=0.76
r184 3 51 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.37 $X2=2.595 $Y2=0.76
r185 2 35 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=1.455
+ $Y=0.37 $X2=1.595 $Y2=0.76
r186 1 85 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_8%VPWR 1 2 3 4 5 6 21 25 29 31 35 39 41 43 47
+ 49 57 62 67 75 81 84 87 90 93 97
r129 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r130 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r131 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r132 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r133 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r134 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r135 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 79 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r137 79 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r138 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r139 76 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=3.33
+ $X2=9.33 $Y2=3.33
r140 76 78 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.495 $Y=3.33
+ $X2=9.84 $Y2=3.33
r141 75 96 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.115 $Y=3.33
+ $X2=10.337 $Y2=3.33
r142 75 78 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=3.33
+ $X2=9.84 $Y2=3.33
r143 74 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r144 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r145 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r146 71 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r147 70 73 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r148 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r149 68 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.735 $Y=3.33
+ $X2=7.57 $Y2=3.33
r150 68 70 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.735 $Y=3.33
+ $X2=7.92 $Y2=3.33
r151 67 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.165 $Y=3.33
+ $X2=9.33 $Y2=3.33
r152 67 73 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.165 $Y=3.33
+ $X2=8.88 $Y2=3.33
r153 66 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r154 66 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r155 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r156 63 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=5.535 $Y2=3.33
r157 63 65 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.7 $Y=3.33 $X2=6
+ $Y2=3.33
r158 62 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.37 $Y=3.33
+ $X2=6.535 $Y2=3.33
r159 62 65 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.37 $Y=3.33 $X2=6
+ $Y2=3.33
r160 61 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r161 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r162 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.7 $Y=3.33
+ $X2=4.535 $Y2=3.33
r163 58 60 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.7 $Y=3.33
+ $X2=5.04 $Y2=3.33
r164 57 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=3.33
+ $X2=5.535 $Y2=3.33
r165 57 60 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.37 $Y=3.33
+ $X2=5.04 $Y2=3.33
r166 56 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r167 55 56 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 52 56 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r169 51 55 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r170 51 52 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r171 49 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.535 $Y2=3.33
r172 49 55 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.08 $Y2=3.33
r173 47 85 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r174 47 61 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r175 43 46 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.28 $Y=2.145
+ $X2=10.28 $Y2=2.825
r176 41 96 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.28 $Y=3.245
+ $X2=10.337 $Y2=3.33
r177 41 46 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=10.28 $Y=3.245
+ $X2=10.28 $Y2=2.825
r178 37 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.33 $Y=3.245
+ $X2=9.33 $Y2=3.33
r179 37 39 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=9.33 $Y=3.245
+ $X2=9.33 $Y2=2.72
r180 33 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.57 $Y=3.245
+ $X2=7.57 $Y2=3.33
r181 33 35 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=7.57 $Y=3.245
+ $X2=7.57 $Y2=2.985
r182 32 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.7 $Y=3.33
+ $X2=6.535 $Y2=3.33
r183 31 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=3.33
+ $X2=7.57 $Y2=3.33
r184 31 32 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.405 $Y=3.33
+ $X2=6.7 $Y2=3.33
r185 27 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.535 $Y=3.245
+ $X2=6.535 $Y2=3.33
r186 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.535 $Y=3.245
+ $X2=6.535 $Y2=2.815
r187 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=3.245
+ $X2=5.535 $Y2=3.33
r188 23 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.535 $Y=3.245
+ $X2=5.535 $Y2=2.815
r189 19 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.535 $Y=3.245
+ $X2=4.535 $Y2=3.33
r190 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.535 $Y=3.245
+ $X2=4.535 $Y2=2.815
r191 6 46 400 $w=1.7e-07 $l=1.05734e-06 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=1.84 $X2=10.28 $Y2=2.825
r192 6 43 400 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=1.84 $X2=10.28 $Y2=2.145
r193 5 39 600 $w=1.7e-07 $l=9.5205e-07 $layer=licon1_PDIFF $count=1 $X=9.18
+ $Y=1.84 $X2=9.33 $Y2=2.72
r194 4 35 600 $w=1.7e-07 $l=1.25702e-06 $layer=licon1_PDIFF $count=1 $X=7.335
+ $Y=1.84 $X2=7.57 $Y2=2.985
r195 3 29 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=6.335
+ $Y=1.84 $X2=6.535 $Y2=2.815
r196 2 25 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.84 $X2=5.535 $Y2=2.815
r197 1 21 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=1.84 $X2=4.535 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_8%A_27_74# 1 2 3 4 5 6 7 8 9 30 32 33 36 38 42
+ 44 48 50 55 56 57 60 62 66 68 72 74 78 80 81 82 83 87 88
c165 83 0 1.96005e-20 $X=4.885 $Y=1.225
c166 56 0 2.61838e-20 $X=4.72 $Y=1.225
r167 83 85 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.885 $Y=1.225
+ $X2=4.885 $Y2=1.385
r168 83 84 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=1.225
+ $X2=4.885 $Y2=1.14
r169 76 78 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=7.425 $Y=1.3
+ $X2=7.425 $Y2=0.515
r170 75 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.69 $Y=1.385
+ $X2=6.565 $Y2=1.385
r171 74 76 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.3 $Y=1.385
+ $X2=7.425 $Y2=1.3
r172 74 75 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.3 $Y=1.385
+ $X2=6.69 $Y2=1.385
r173 70 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.565 $Y=1.3
+ $X2=6.565 $Y2=1.385
r174 70 72 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=6.565 $Y=1.3
+ $X2=6.565 $Y2=0.515
r175 69 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.83 $Y=1.385
+ $X2=5.705 $Y2=1.385
r176 68 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.44 $Y=1.385
+ $X2=6.565 $Y2=1.385
r177 68 69 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.44 $Y=1.385
+ $X2=5.83 $Y2=1.385
r178 64 87 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.705 $Y=1.3
+ $X2=5.705 $Y2=1.385
r179 64 66 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=5.705 $Y=1.3
+ $X2=5.705 $Y2=0.515
r180 63 85 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.05 $Y=1.385
+ $X2=4.885 $Y2=1.385
r181 62 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.58 $Y=1.385
+ $X2=5.705 $Y2=1.385
r182 62 63 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.58 $Y=1.385
+ $X2=5.05 $Y2=1.385
r183 60 84 28.8111 $w=2.48e-07 $l=6.25e-07 $layer=LI1_cond $X=4.925 $Y=0.515
+ $X2=4.925 $Y2=1.14
r184 56 83 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.72 $Y=1.225
+ $X2=4.885 $Y2=1.225
r185 56 57 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.72 $Y=1.225
+ $X2=4.11 $Y2=1.225
r186 53 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.025 $Y=1.14
+ $X2=4.11 $Y2=1.225
r187 53 55 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.025 $Y=1.14
+ $X2=4.025 $Y2=0.515
r188 52 55 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.025 $Y=0.425
+ $X2=4.025 $Y2=0.515
r189 51 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=0.34
+ $X2=3.095 $Y2=0.34
r190 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.94 $Y=0.34
+ $X2=4.025 $Y2=0.425
r191 50 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.94 $Y=0.34
+ $X2=3.26 $Y2=0.34
r192 46 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.425
+ $X2=3.095 $Y2=0.34
r193 46 48 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.095 $Y=0.425
+ $X2=3.095 $Y2=0.645
r194 45 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0.34
+ $X2=2.095 $Y2=0.34
r195 44 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=0.34
+ $X2=3.095 $Y2=0.34
r196 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.93 $Y=0.34
+ $X2=2.26 $Y2=0.34
r197 40 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.425
+ $X2=2.095 $Y2=0.34
r198 40 42 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.095 $Y=0.425
+ $X2=2.095 $Y2=0.645
r199 39 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.34
+ $X2=1.14 $Y2=0.34
r200 38 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=0.34
+ $X2=2.095 $Y2=0.34
r201 38 39 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.93 $Y=0.34
+ $X2=1.225 $Y2=0.34
r202 34 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.425
+ $X2=1.14 $Y2=0.34
r203 34 36 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.14 $Y=0.425
+ $X2=1.14 $Y2=0.63
r204 32 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=0.34
+ $X2=1.14 $Y2=0.34
r205 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=0.34
+ $X2=0.365 $Y2=0.34
r206 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.365 $Y2=0.34
r207 28 30 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.24 $Y2=0.515
r208 9 78 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.325
+ $Y=0.37 $X2=7.465 $Y2=0.515
r209 8 72 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.465
+ $Y=0.37 $X2=6.605 $Y2=0.515
r210 7 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.605
+ $Y=0.37 $X2=5.745 $Y2=0.515
r211 6 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.745
+ $Y=0.37 $X2=4.885 $Y2=0.515
r212 5 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.37 $X2=4.025 $Y2=0.515
r213 4 48 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=2.885
+ $Y=0.37 $X2=3.095 $Y2=0.645
r214 3 42 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=1.885
+ $Y=0.37 $X2=2.095 $Y2=0.645
r215 2 36 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.63
r216 1 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_8%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 47 48 50 51 52 67 71 76 82 85 89
c130 21 0 1.9142e-19 $X=4.455 $Y=0.495
r131 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r132 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r133 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r134 80 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r135 80 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r136 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r137 77 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.5 $Y=0 $X2=9.415
+ $Y2=0
r138 77 79 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.5 $Y=0 $X2=9.84
+ $Y2=0
r139 76 88 4.77426 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=10.11 $Y=0
+ $X2=10.335 $Y2=0
r140 76 79 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=10.11 $Y=0 $X2=9.84
+ $Y2=0
r141 75 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=9.36 $Y2=0
r142 75 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r143 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r144 72 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.12 $Y=0 $X2=6.995
+ $Y2=0
r145 72 74 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.12 $Y=0 $X2=7.44
+ $Y2=0
r146 71 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.33 $Y=0 $X2=9.415
+ $Y2=0
r147 71 74 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=9.33 $Y=0 $X2=7.44
+ $Y2=0
r148 70 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r149 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r150 67 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.87 $Y=0 $X2=6.995
+ $Y2=0
r151 67 69 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.87 $Y=0 $X2=6.48
+ $Y2=0
r152 66 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r153 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r154 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r155 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r156 59 60 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r157 56 60 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r158 55 59 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r159 55 56 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r160 52 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=6
+ $Y2=0
r161 52 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.04 $Y2=0
r162 50 65 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.01 $Y=0 $X2=6
+ $Y2=0
r163 50 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.01 $Y=0 $X2=6.135
+ $Y2=0
r164 49 69 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.26 $Y=0 $X2=6.48
+ $Y2=0
r165 49 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.26 $Y=0 $X2=6.135
+ $Y2=0
r166 47 62 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.04
+ $Y2=0
r167 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.315
+ $Y2=0
r168 46 65 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.4 $Y=0 $X2=6 $Y2=0
r169 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=0 $X2=5.315
+ $Y2=0
r170 44 59 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.08
+ $Y2=0
r171 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.455
+ $Y2=0
r172 43 62 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.62 $Y=0 $X2=5.04
+ $Y2=0
r173 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=0 $X2=4.455
+ $Y2=0
r174 39 88 3.03431 $w=3.35e-07 $l=1.1025e-07 $layer=LI1_cond $X=10.277 $Y=0.085
+ $X2=10.335 $Y2=0
r175 39 41 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=10.277 $Y=0.085
+ $X2=10.277 $Y2=0.515
r176 35 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.415 $Y=0.085
+ $X2=9.415 $Y2=0
r177 35 37 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.415 $Y=0.085
+ $X2=9.415 $Y2=0.505
r178 31 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=0.085
+ $X2=6.995 $Y2=0
r179 31 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.995 $Y=0.085
+ $X2=6.995 $Y2=0.515
r180 27 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.135 $Y=0.085
+ $X2=6.135 $Y2=0
r181 27 29 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.135 $Y=0.085
+ $X2=6.135 $Y2=0.515
r182 23 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=0.085
+ $X2=5.315 $Y2=0
r183 23 25 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.315 $Y=0.085
+ $X2=5.315 $Y2=0.515
r184 19 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0.085
+ $X2=4.455 $Y2=0
r185 19 21 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.455 $Y=0.085
+ $X2=4.455 $Y2=0.495
r186 6 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=10.135
+ $Y=0.37 $X2=10.275 $Y2=0.515
r187 5 37 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=9.275
+ $Y=0.37 $X2=9.415 $Y2=0.505
r188 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.895
+ $Y=0.37 $X2=7.035 $Y2=0.515
r189 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.035
+ $Y=0.37 $X2=6.175 $Y2=0.515
r190 2 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.175
+ $Y=0.37 $X2=5.315 $Y2=0.515
r191 1 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.315
+ $Y=0.37 $X2=4.455 $Y2=0.495
.ends

