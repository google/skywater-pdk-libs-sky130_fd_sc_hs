* File: sky130_fd_sc_hs__and2_4.pxi.spice
* Created: Thu Aug 27 20:31:46 2020
* 
x_PM_SKY130_FD_SC_HS__AND2_4%A_83_269# N_A_83_269#_M1005_d N_A_83_269#_M1000_d
+ N_A_83_269#_M1007_d N_A_83_269#_c_84_n N_A_83_269#_M1002_g N_A_83_269#_c_94_n
+ N_A_83_269#_M1003_g N_A_83_269#_c_85_n N_A_83_269#_M1004_g N_A_83_269#_c_95_n
+ N_A_83_269#_M1012_g N_A_83_269#_c_86_n N_A_83_269#_M1008_g N_A_83_269#_c_96_n
+ N_A_83_269#_M1013_g N_A_83_269#_c_97_n N_A_83_269#_M1014_g N_A_83_269#_c_87_n
+ N_A_83_269#_M1015_g N_A_83_269#_c_88_n N_A_83_269#_c_98_n N_A_83_269#_c_99_n
+ N_A_83_269#_c_147_p N_A_83_269#_c_100_n N_A_83_269#_c_101_n N_A_83_269#_c_89_n
+ N_A_83_269#_c_90_n N_A_83_269#_c_91_n N_A_83_269#_c_92_n N_A_83_269#_c_103_n
+ N_A_83_269#_c_104_n N_A_83_269#_c_105_n N_A_83_269#_c_93_n
+ PM_SKY130_FD_SC_HS__AND2_4%A_83_269#
x_PM_SKY130_FD_SC_HS__AND2_4%A N_A_c_235_n N_A_M1001_g N_A_M1005_g N_A_c_236_n
+ N_A_M1007_g N_A_M1010_g A N_A_c_234_n PM_SKY130_FD_SC_HS__AND2_4%A
x_PM_SKY130_FD_SC_HS__AND2_4%B N_B_c_287_n N_B_c_288_n N_B_M1000_g N_B_M1009_g
+ N_B_c_280_n N_B_c_281_n N_B_c_282_n N_B_c_283_n N_B_c_290_n N_B_M1006_g
+ N_B_M1011_g B N_B_c_286_n PM_SKY130_FD_SC_HS__AND2_4%B
x_PM_SKY130_FD_SC_HS__AND2_4%VPWR N_VPWR_M1003_d N_VPWR_M1012_d N_VPWR_M1014_d
+ N_VPWR_M1001_s N_VPWR_M1006_s N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n
+ N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_362_n
+ N_VPWR_c_363_n VPWR N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n
+ N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_354_n PM_SKY130_FD_SC_HS__AND2_4%VPWR
x_PM_SKY130_FD_SC_HS__AND2_4%X N_X_M1002_s N_X_M1008_s N_X_M1003_s N_X_M1013_s
+ N_X_c_427_n N_X_c_430_n N_X_c_437_n N_X_c_442_n N_X_c_446_n N_X_c_431_n
+ N_X_c_428_n N_X_c_457_n N_X_c_458_n X N_X_c_429_n X
+ PM_SKY130_FD_SC_HS__AND2_4%X
x_PM_SKY130_FD_SC_HS__AND2_4%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_M1015_d
+ N_VGND_M1011_s N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n N_VGND_c_494_n
+ N_VGND_c_495_n N_VGND_c_496_n VGND N_VGND_c_497_n N_VGND_c_498_n
+ N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n
+ PM_SKY130_FD_SC_HS__AND2_4%VGND
x_PM_SKY130_FD_SC_HS__AND2_4%A_504_119# N_A_504_119#_M1009_d
+ N_A_504_119#_M1010_s N_A_504_119#_c_551_n N_A_504_119#_c_552_n
+ N_A_504_119#_c_553_n N_A_504_119#_c_554_n
+ PM_SKY130_FD_SC_HS__AND2_4%A_504_119#
cc_1 VNB N_A_83_269#_c_84_n 0.0190055f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_2 VNB N_A_83_269#_c_85_n 0.0157541f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.345
cc_3 VNB N_A_83_269#_c_86_n 0.0171136f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.345
cc_4 VNB N_A_83_269#_c_87_n 0.0180145f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.345
cc_5 VNB N_A_83_269#_c_88_n 0.00247544f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=1.51
cc_6 VNB N_A_83_269#_c_89_n 0.0012516f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=0.72
cc_7 VNB N_A_83_269#_c_90_n 0.00120857f $X=-0.19 $Y=-0.245 $X2=3.5 $Y2=1.195
cc_8 VNB N_A_83_269#_c_91_n 0.00327749f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=1.195
cc_9 VNB N_A_83_269#_c_92_n 0.00784369f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.95
cc_10 VNB N_A_83_269#_c_93_n 0.0874615f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.555
cc_11 VNB N_A_M1005_g 0.0211437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1010_g 0.0206639f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_13 VNB A 0.00134224f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_14 VNB N_A_c_234_n 0.0271196f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.345
cc_15 VNB N_B_M1009_g 0.0267987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_280_n 0.096137f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_17 VNB N_B_c_281_n 0.012503f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.865
cc_18 VNB N_B_c_282_n 0.00935751f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.865
cc_19 VNB N_B_c_283_n 0.0221782f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_20 VNB N_B_M1011_g 0.0277901f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_21 VNB B 0.00598581f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.345
cc_22 VNB N_B_c_286_n 0.02407f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.765
cc_23 VNB N_VPWR_c_354_n 0.183584f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.555
cc_24 VNB N_X_c_427_n 0.00250594f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_25 VNB N_X_c_428_n 0.00304013f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.865
cc_26 VNB N_X_c_429_n 0.00103798f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=2.19
cc_27 VNB N_VGND_c_491_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_28 VNB N_VGND_c_492_n 0.0510645f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_29 VNB N_VGND_c_493_n 0.0108434f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_30 VNB N_VGND_c_494_n 0.0133746f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.865
cc_31 VNB N_VGND_c_495_n 0.0110036f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.765
cc_32 VNB N_VGND_c_496_n 0.0551896f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_33 VNB N_VGND_c_497_n 0.0178324f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.345
cc_34 VNB N_VGND_c_498_n 0.02006f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.51
cc_35 VNB N_VGND_c_499_n 0.0373297f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.51
cc_36 VNB N_VGND_c_500_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=0.72
cc_37 VNB N_VGND_c_501_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.5 $Y2=1.195
cc_38 VNB N_VGND_c_502_n 0.256254f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=2.12
cc_39 VNB N_A_504_119#_c_551_n 0.00348835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_504_119#_c_552_n 0.0172345f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.865
cc_41 VNB N_A_504_119#_c_553_n 7.85965e-19 $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.865
cc_42 VNB N_A_504_119#_c_554_n 0.00459367f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_43 VPB N_A_83_269#_c_94_n 0.0174275f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_44 VPB N_A_83_269#_c_95_n 0.0150815f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_45 VPB N_A_83_269#_c_96_n 0.0157677f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_46 VPB N_A_83_269#_c_97_n 0.0163792f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.765
cc_47 VPB N_A_83_269#_c_98_n 0.00131251f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.95
cc_48 VPB N_A_83_269#_c_99_n 0.00178628f $X=-0.19 $Y=1.66 $X2=2.47 $Y2=2.035
cc_49 VPB N_A_83_269#_c_100_n 0.003262f $X=-0.19 $Y=1.66 $X2=2.635 $Y2=2.19
cc_50 VPB N_A_83_269#_c_101_n 0.00248957f $X=-0.19 $Y=1.66 $X2=3.5 $Y2=2.035
cc_51 VPB N_A_83_269#_c_92_n 0.00588088f $X=-0.19 $Y=1.66 $X2=3.585 $Y2=1.95
cc_52 VPB N_A_83_269#_c_103_n 0.00200197f $X=-0.19 $Y=1.66 $X2=3.585 $Y2=2.19
cc_53 VPB N_A_83_269#_c_104_n 0.00377621f $X=-0.19 $Y=1.66 $X2=2.635 $Y2=2.035
cc_54 VPB N_A_83_269#_c_105_n 0.0010739f $X=-0.19 $Y=1.66 $X2=3.585 $Y2=2.035
cc_55 VPB N_A_83_269#_c_93_n 0.0540219f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.555
cc_56 VPB N_A_c_235_n 0.0146537f $X=-0.19 $Y=1.66 $X2=2.975 $Y2=0.595
cc_57 VPB N_A_c_236_n 0.0139488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_c_234_n 0.0424369f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.345
cc_59 VPB N_B_c_287_n 0.011191f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.045
cc_60 VPB N_B_c_288_n 0.0212431f $X=-0.19 $Y=1.66 $X2=3.435 $Y2=2.045
cc_61 VPB N_B_c_283_n 0.018753f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_62 VPB N_B_c_290_n 0.027016f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_63 VPB B 0.00449364f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.345
cc_64 VPB N_B_c_286_n 0.00513926f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_65 VPB N_VPWR_c_355_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.345
cc_66 VPB N_VPWR_c_356_n 0.057703f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.865
cc_67 VPB N_VPWR_c_357_n 0.0044818f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.865
cc_68 VPB N_VPWR_c_358_n 0.00876009f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.765
cc_69 VPB N_VPWR_c_359_n 0.0102828f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=1.51
cc_70 VPB N_VPWR_c_360_n 0.0123504f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.51
cc_71 VPB N_VPWR_c_361_n 0.0590218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_362_n 0.0183691f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=1.51
cc_73 VPB N_VPWR_c_363_n 0.00460249f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.675
cc_74 VPB N_VPWR_c_364_n 0.0191617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_365_n 0.0201594f $X=-0.19 $Y=1.66 $X2=3.16 $Y2=0.72
cc_76 VPB N_VPWR_c_366_n 0.0169422f $X=-0.19 $Y=1.66 $X2=3.585 $Y2=1.28
cc_77 VPB N_VPWR_c_367_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.555
cc_78 VPB N_VPWR_c_368_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.555
cc_79 VPB N_VPWR_c_354_n 0.0831938f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.555
cc_80 VPB N_X_c_430_n 0.00217015f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_81 VPB N_X_c_431_n 0.00217444f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=2.4
cc_82 VPB X 0.00138178f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.675
cc_83 N_A_83_269#_c_100_n N_A_c_235_n 0.00101488f $X=2.635 $Y=2.19 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_83_269#_c_101_n N_A_c_235_n 0.011583f $X=3.5 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_83_269#_c_91_n N_A_M1005_g 0.00146831f $X=3.325 $Y=1.195 $X2=0 $Y2=0
cc_86 N_A_83_269#_c_101_n N_A_c_236_n 0.0109536f $X=3.5 $Y=2.035 $X2=0 $Y2=0
cc_87 N_A_83_269#_c_103_n N_A_c_236_n 0.00601403f $X=3.585 $Y=2.19 $X2=0 $Y2=0
cc_88 N_A_83_269#_c_89_n N_A_M1010_g 0.00677769f $X=3.16 $Y=0.72 $X2=0 $Y2=0
cc_89 N_A_83_269#_c_90_n N_A_M1010_g 0.0123722f $X=3.5 $Y=1.195 $X2=0 $Y2=0
cc_90 N_A_83_269#_c_91_n N_A_M1010_g 0.00157603f $X=3.325 $Y=1.195 $X2=0 $Y2=0
cc_91 N_A_83_269#_c_92_n N_A_M1010_g 0.0115076f $X=3.585 $Y=1.95 $X2=0 $Y2=0
cc_92 N_A_83_269#_c_101_n A 0.0245865f $X=3.5 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_83_269#_c_91_n A 0.0219645f $X=3.325 $Y=1.195 $X2=0 $Y2=0
cc_94 N_A_83_269#_c_92_n A 0.0188613f $X=3.585 $Y=1.95 $X2=0 $Y2=0
cc_95 N_A_83_269#_c_101_n N_A_c_234_n 0.0222872f $X=3.5 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_83_269#_c_91_n N_A_c_234_n 0.00113662f $X=3.325 $Y=1.195 $X2=0 $Y2=0
cc_97 N_A_83_269#_c_104_n N_A_c_234_n 6.13048e-19 $X=2.635 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_83_269#_c_97_n N_B_c_287_n 0.00591137f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_83_269#_c_98_n N_B_c_287_n 0.00359939f $X=1.97 $Y=1.95 $X2=0 $Y2=0
cc_100 N_A_83_269#_c_93_n N_B_c_287_n 0.002946f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_101 N_A_83_269#_c_97_n N_B_c_288_n 0.017545f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_83_269#_c_99_n N_B_c_288_n 0.0128428f $X=2.47 $Y=2.035 $X2=0 $Y2=0
cc_103 N_A_83_269#_c_100_n N_B_c_288_n 0.0118949f $X=2.635 $Y=2.19 $X2=0 $Y2=0
cc_104 N_A_83_269#_c_104_n N_B_c_288_n 0.00227727f $X=2.635 $Y=2.035 $X2=0 $Y2=0
cc_105 N_A_83_269#_c_87_n N_B_M1009_g 0.0176506f $X=1.935 $Y=1.345 $X2=0 $Y2=0
cc_106 N_A_83_269#_c_92_n N_B_c_282_n 0.0153689f $X=3.585 $Y=1.95 $X2=0 $Y2=0
cc_107 N_A_83_269#_c_103_n N_B_c_290_n 0.00326147f $X=3.585 $Y=2.19 $X2=0 $Y2=0
cc_108 N_A_83_269#_c_105_n N_B_c_290_n 0.00287096f $X=3.585 $Y=2.035 $X2=0 $Y2=0
cc_109 N_A_83_269#_c_89_n N_B_M1011_g 5.82683e-19 $X=3.16 $Y=0.72 $X2=0 $Y2=0
cc_110 N_A_83_269#_c_90_n N_B_M1011_g 0.00200207f $X=3.5 $Y=1.195 $X2=0 $Y2=0
cc_111 N_A_83_269#_c_92_n N_B_M1011_g 6.77794e-19 $X=3.585 $Y=1.95 $X2=0 $Y2=0
cc_112 N_A_83_269#_c_88_n B 0.0253761f $X=1.885 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A_83_269#_c_98_n B 0.0076003f $X=1.97 $Y=1.95 $X2=0 $Y2=0
cc_114 N_A_83_269#_c_99_n B 0.0161894f $X=2.47 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A_83_269#_c_104_n B 0.0254551f $X=2.635 $Y=2.035 $X2=0 $Y2=0
cc_116 N_A_83_269#_c_93_n B 6.88662e-19 $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_117 N_A_83_269#_c_88_n N_B_c_286_n 0.00133751f $X=1.885 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A_83_269#_c_99_n N_B_c_286_n 3.50421e-19 $X=2.47 $Y=2.035 $X2=0 $Y2=0
cc_119 N_A_83_269#_c_104_n N_B_c_286_n 5.16717e-19 $X=2.635 $Y=2.035 $X2=0 $Y2=0
cc_120 N_A_83_269#_c_93_n N_B_c_286_n 0.0182298f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_121 N_A_83_269#_c_98_n N_VPWR_M1014_d 0.00135982f $X=1.97 $Y=1.95 $X2=0 $Y2=0
cc_122 N_A_83_269#_c_99_n N_VPWR_M1014_d 0.00890498f $X=2.47 $Y=2.035 $X2=0
+ $Y2=0
cc_123 N_A_83_269#_c_147_p N_VPWR_M1014_d 5.20113e-19 $X=2.055 $Y=2.035 $X2=0
+ $Y2=0
cc_124 N_A_83_269#_c_101_n N_VPWR_M1001_s 0.00224297f $X=3.5 $Y=2.035 $X2=0
+ $Y2=0
cc_125 N_A_83_269#_c_94_n N_VPWR_c_356_n 0.00841517f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_83_269#_c_94_n N_VPWR_c_357_n 6.00285e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A_83_269#_c_95_n N_VPWR_c_357_n 0.0125784f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A_83_269#_c_96_n N_VPWR_c_357_n 0.00466682f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A_83_269#_c_96_n N_VPWR_c_358_n 5.72968e-19 $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_83_269#_c_97_n N_VPWR_c_358_n 0.0121347f $X=1.875 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_83_269#_c_99_n N_VPWR_c_358_n 0.0169675f $X=2.47 $Y=2.035 $X2=0 $Y2=0
cc_132 N_A_83_269#_c_147_p N_VPWR_c_358_n 0.00542547f $X=2.055 $Y=2.035 $X2=0
+ $Y2=0
cc_133 N_A_83_269#_c_100_n N_VPWR_c_358_n 0.0413658f $X=2.635 $Y=2.19 $X2=0
+ $Y2=0
cc_134 N_A_83_269#_c_100_n N_VPWR_c_359_n 0.00158095f $X=2.635 $Y=2.19 $X2=0
+ $Y2=0
cc_135 N_A_83_269#_c_101_n N_VPWR_c_359_n 0.0181909f $X=3.5 $Y=2.035 $X2=0 $Y2=0
cc_136 N_A_83_269#_c_103_n N_VPWR_c_359_n 0.0400865f $X=3.585 $Y=2.19 $X2=0
+ $Y2=0
cc_137 N_A_83_269#_c_103_n N_VPWR_c_361_n 0.0511276f $X=3.585 $Y=2.19 $X2=0
+ $Y2=0
cc_138 N_A_83_269#_c_105_n N_VPWR_c_361_n 0.00695516f $X=3.585 $Y=2.035 $X2=0
+ $Y2=0
cc_139 N_A_83_269#_c_94_n N_VPWR_c_362_n 0.00422942f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_83_269#_c_95_n N_VPWR_c_362_n 0.00413917f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A_83_269#_c_96_n N_VPWR_c_364_n 0.00445602f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_83_269#_c_97_n N_VPWR_c_364_n 0.00413917f $X=1.875 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_83_269#_c_100_n N_VPWR_c_365_n 0.0111926f $X=2.635 $Y=2.19 $X2=0
+ $Y2=0
cc_144 N_A_83_269#_c_103_n N_VPWR_c_366_n 0.00575213f $X=3.585 $Y=2.19 $X2=0
+ $Y2=0
cc_145 N_A_83_269#_c_94_n N_VPWR_c_354_n 0.0078771f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_83_269#_c_95_n N_VPWR_c_354_n 0.00817726f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_83_269#_c_96_n N_VPWR_c_354_n 0.00857779f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_83_269#_c_97_n N_VPWR_c_354_n 0.00817916f $X=1.875 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_A_83_269#_c_100_n N_VPWR_c_354_n 0.0115381f $X=2.635 $Y=2.19 $X2=0
+ $Y2=0
cc_150 N_A_83_269#_c_103_n N_VPWR_c_354_n 0.00591657f $X=3.585 $Y=2.19 $X2=0
+ $Y2=0
cc_151 N_A_83_269#_c_84_n N_X_c_427_n 0.0068035f $X=0.495 $Y=1.345 $X2=0 $Y2=0
cc_152 N_A_83_269#_c_85_n N_X_c_427_n 3.97481e-19 $X=0.925 $Y=1.345 $X2=0 $Y2=0
cc_153 N_A_83_269#_c_94_n N_X_c_430_n 0.0119433f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_83_269#_c_95_n N_X_c_430_n 0.0045777f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_83_269#_c_85_n N_X_c_437_n 0.014204f $X=0.925 $Y=1.345 $X2=0 $Y2=0
cc_156 N_A_83_269#_c_86_n N_X_c_437_n 0.0143843f $X=1.355 $Y=1.345 $X2=0 $Y2=0
cc_157 N_A_83_269#_c_87_n N_X_c_437_n 0.00170179f $X=1.935 $Y=1.345 $X2=0 $Y2=0
cc_158 N_A_83_269#_c_88_n N_X_c_437_n 0.0488551f $X=1.885 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A_83_269#_c_93_n N_X_c_437_n 0.00701064f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_160 N_A_83_269#_c_95_n N_X_c_442_n 0.0144622f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_83_269#_c_96_n N_X_c_442_n 0.0120074f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_83_269#_c_88_n N_X_c_442_n 0.0294034f $X=1.885 $Y=1.51 $X2=0 $Y2=0
cc_163 N_A_83_269#_c_93_n N_X_c_442_n 0.00653905f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_164 N_A_83_269#_c_96_n N_X_c_446_n 3.69071e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_83_269#_c_88_n N_X_c_446_n 0.0180035f $X=1.885 $Y=1.51 $X2=0 $Y2=0
cc_166 N_A_83_269#_c_98_n N_X_c_446_n 0.00825359f $X=1.97 $Y=1.95 $X2=0 $Y2=0
cc_167 N_A_83_269#_c_147_p N_X_c_446_n 0.00568121f $X=2.055 $Y=2.035 $X2=0 $Y2=0
cc_168 N_A_83_269#_c_93_n N_X_c_446_n 0.00509567f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_169 N_A_83_269#_c_95_n N_X_c_431_n 7.37455e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A_83_269#_c_96_n N_X_c_431_n 0.0118193f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_83_269#_c_97_n N_X_c_431_n 0.00651572f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_83_269#_c_147_p N_X_c_431_n 0.00844191f $X=2.055 $Y=2.035 $X2=0 $Y2=0
cc_173 N_A_83_269#_c_86_n N_X_c_428_n 0.00334069f $X=1.355 $Y=1.345 $X2=0 $Y2=0
cc_174 N_A_83_269#_c_87_n N_X_c_428_n 0.00474848f $X=1.935 $Y=1.345 $X2=0 $Y2=0
cc_175 N_A_83_269#_c_84_n N_X_c_457_n 0.00186215f $X=0.495 $Y=1.345 $X2=0 $Y2=0
cc_176 N_A_83_269#_c_94_n N_X_c_458_n 0.00197815f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_83_269#_c_94_n X 0.00337225f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_83_269#_c_95_n X 0.0020009f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A_83_269#_c_88_n X 0.00980665f $X=1.885 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_83_269#_c_93_n X 0.0244979f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_181 N_A_83_269#_c_84_n N_X_c_429_n 0.00559035f $X=0.495 $Y=1.345 $X2=0 $Y2=0
cc_182 N_A_83_269#_c_85_n N_X_c_429_n 0.00280039f $X=0.925 $Y=1.345 $X2=0 $Y2=0
cc_183 N_A_83_269#_c_88_n N_X_c_429_n 0.0134383f $X=1.885 $Y=1.51 $X2=0 $Y2=0
cc_184 N_A_83_269#_c_93_n N_X_c_429_n 0.0185187f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_185 N_A_83_269#_c_84_n N_VGND_c_492_n 0.00513328f $X=0.495 $Y=1.345 $X2=0
+ $Y2=0
cc_186 N_A_83_269#_c_84_n N_VGND_c_493_n 4.50936e-19 $X=0.495 $Y=1.345 $X2=0
+ $Y2=0
cc_187 N_A_83_269#_c_85_n N_VGND_c_493_n 0.00819261f $X=0.925 $Y=1.345 $X2=0
+ $Y2=0
cc_188 N_A_83_269#_c_86_n N_VGND_c_493_n 0.00838873f $X=1.355 $Y=1.345 $X2=0
+ $Y2=0
cc_189 N_A_83_269#_c_87_n N_VGND_c_493_n 5.69258e-19 $X=1.935 $Y=1.345 $X2=0
+ $Y2=0
cc_190 N_A_83_269#_c_86_n N_VGND_c_494_n 7.80783e-19 $X=1.355 $Y=1.345 $X2=0
+ $Y2=0
cc_191 N_A_83_269#_c_87_n N_VGND_c_494_n 0.0135521f $X=1.935 $Y=1.345 $X2=0
+ $Y2=0
cc_192 N_A_83_269#_c_88_n N_VGND_c_494_n 0.00407487f $X=1.885 $Y=1.51 $X2=0
+ $Y2=0
cc_193 N_A_83_269#_c_89_n N_VGND_c_496_n 0.00484906f $X=3.16 $Y=0.72 $X2=0 $Y2=0
cc_194 N_A_83_269#_c_90_n N_VGND_c_496_n 0.0103921f $X=3.5 $Y=1.195 $X2=0 $Y2=0
cc_195 N_A_83_269#_c_84_n N_VGND_c_497_n 0.00470409f $X=0.495 $Y=1.345 $X2=0
+ $Y2=0
cc_196 N_A_83_269#_c_85_n N_VGND_c_497_n 0.00407914f $X=0.925 $Y=1.345 $X2=0
+ $Y2=0
cc_197 N_A_83_269#_c_86_n N_VGND_c_498_n 0.00407914f $X=1.355 $Y=1.345 $X2=0
+ $Y2=0
cc_198 N_A_83_269#_c_87_n N_VGND_c_498_n 0.00407914f $X=1.935 $Y=1.345 $X2=0
+ $Y2=0
cc_199 N_A_83_269#_c_84_n N_VGND_c_502_n 0.00506877f $X=0.495 $Y=1.345 $X2=0
+ $Y2=0
cc_200 N_A_83_269#_c_85_n N_VGND_c_502_n 0.00425776f $X=0.925 $Y=1.345 $X2=0
+ $Y2=0
cc_201 N_A_83_269#_c_86_n N_VGND_c_502_n 0.00425776f $X=1.355 $Y=1.345 $X2=0
+ $Y2=0
cc_202 N_A_83_269#_c_87_n N_VGND_c_502_n 0.00425776f $X=1.935 $Y=1.345 $X2=0
+ $Y2=0
cc_203 N_A_83_269#_c_90_n N_A_504_119#_M1010_s 0.00322345f $X=3.5 $Y=1.195 $X2=0
+ $Y2=0
cc_204 N_A_83_269#_c_87_n N_A_504_119#_c_551_n 2.18891e-19 $X=1.935 $Y=1.345
+ $X2=0 $Y2=0
cc_205 N_A_83_269#_c_89_n N_A_504_119#_c_552_n 0.0216292f $X=3.16 $Y=0.72 $X2=0
+ $Y2=0
cc_206 N_A_83_269#_c_90_n N_A_504_119#_c_554_n 0.0147044f $X=3.5 $Y=1.195 $X2=0
+ $Y2=0
cc_207 N_A_c_234_n N_B_c_287_n 0.0143436f $X=3.36 $Y=1.71 $X2=0 $Y2=0
cc_208 N_A_c_235_n N_B_c_288_n 0.012455f $X=2.885 $Y=1.97 $X2=0 $Y2=0
cc_209 N_A_M1005_g N_B_M1009_g 0.00953605f $X=2.9 $Y=0.915 $X2=0 $Y2=0
cc_210 N_A_M1005_g N_B_c_280_n 0.00882199f $X=2.9 $Y=0.915 $X2=0 $Y2=0
cc_211 N_A_M1010_g N_B_c_280_n 0.00882199f $X=3.375 $Y=0.915 $X2=0 $Y2=0
cc_212 N_A_M1010_g N_B_c_282_n 0.0134112f $X=3.375 $Y=0.915 $X2=0 $Y2=0
cc_213 N_A_c_234_n N_B_c_283_n 0.0134112f $X=3.36 $Y=1.71 $X2=0 $Y2=0
cc_214 N_A_c_236_n N_B_c_290_n 0.0125221f $X=3.36 $Y=1.97 $X2=0 $Y2=0
cc_215 N_A_M1010_g N_B_M1011_g 0.0172255f $X=3.375 $Y=0.915 $X2=0 $Y2=0
cc_216 N_A_M1005_g B 0.00294883f $X=2.9 $Y=0.915 $X2=0 $Y2=0
cc_217 A B 0.0270483f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_218 N_A_c_234_n B 0.00292892f $X=3.36 $Y=1.71 $X2=0 $Y2=0
cc_219 N_A_M1005_g N_B_c_286_n 0.00516243f $X=2.9 $Y=0.915 $X2=0 $Y2=0
cc_220 N_A_c_234_n N_B_c_286_n 0.0145976f $X=3.36 $Y=1.71 $X2=0 $Y2=0
cc_221 N_A_c_235_n N_VPWR_c_359_n 0.00339887f $X=2.885 $Y=1.97 $X2=0 $Y2=0
cc_222 N_A_c_236_n N_VPWR_c_359_n 0.0101707f $X=3.36 $Y=1.97 $X2=0 $Y2=0
cc_223 N_A_c_236_n N_VPWR_c_361_n 6.01201e-19 $X=3.36 $Y=1.97 $X2=0 $Y2=0
cc_224 N_A_c_235_n N_VPWR_c_365_n 0.00523993f $X=2.885 $Y=1.97 $X2=0 $Y2=0
cc_225 N_A_c_236_n N_VPWR_c_366_n 0.00470366f $X=3.36 $Y=1.97 $X2=0 $Y2=0
cc_226 N_A_c_235_n N_VPWR_c_354_n 0.0052212f $X=2.885 $Y=1.97 $X2=0 $Y2=0
cc_227 N_A_c_236_n N_VPWR_c_354_n 0.00473388f $X=3.36 $Y=1.97 $X2=0 $Y2=0
cc_228 N_A_M1010_g N_VGND_c_496_n 7.48424e-19 $X=3.375 $Y=0.915 $X2=0 $Y2=0
cc_229 N_A_M1005_g N_A_504_119#_c_551_n 0.00379535f $X=2.9 $Y=0.915 $X2=0 $Y2=0
cc_230 N_A_M1005_g N_A_504_119#_c_552_n 0.00369782f $X=2.9 $Y=0.915 $X2=0 $Y2=0
cc_231 N_A_M1010_g N_A_504_119#_c_552_n 0.00330666f $X=3.375 $Y=0.915 $X2=0
+ $Y2=0
cc_232 N_A_M1010_g N_A_504_119#_c_554_n 0.00311697f $X=3.375 $Y=0.915 $X2=0
+ $Y2=0
cc_233 N_B_c_288_n N_VPWR_c_358_n 0.00865871f $X=2.41 $Y=1.97 $X2=0 $Y2=0
cc_234 N_B_c_290_n N_VPWR_c_359_n 5.11845e-19 $X=3.81 $Y=1.97 $X2=0 $Y2=0
cc_235 N_B_c_290_n N_VPWR_c_361_n 0.0189904f $X=3.81 $Y=1.97 $X2=0 $Y2=0
cc_236 N_B_c_288_n N_VPWR_c_365_n 0.00510653f $X=2.41 $Y=1.97 $X2=0 $Y2=0
cc_237 N_B_c_290_n N_VPWR_c_366_n 0.00470366f $X=3.81 $Y=1.97 $X2=0 $Y2=0
cc_238 N_B_c_288_n N_VPWR_c_354_n 0.0052212f $X=2.41 $Y=1.97 $X2=0 $Y2=0
cc_239 N_B_c_290_n N_VPWR_c_354_n 0.00473388f $X=3.81 $Y=1.97 $X2=0 $Y2=0
cc_240 N_B_c_281_n N_VGND_c_494_n 0.0133187f $X=2.52 $Y=0.18 $X2=0 $Y2=0
cc_241 B N_VGND_c_494_n 0.0049234f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B_c_286_n N_VGND_c_494_n 0.0013714f $X=2.42 $Y=1.51 $X2=0 $Y2=0
cc_243 N_B_c_280_n N_VGND_c_496_n 0.00763335f $X=3.75 $Y=0.18 $X2=0 $Y2=0
cc_244 N_B_M1011_g N_VGND_c_496_n 0.0206326f $X=3.825 $Y=0.915 $X2=0 $Y2=0
cc_245 N_B_c_281_n N_VGND_c_499_n 0.0368558f $X=2.52 $Y=0.18 $X2=0 $Y2=0
cc_246 N_B_c_280_n N_VGND_c_502_n 0.0391084f $X=3.75 $Y=0.18 $X2=0 $Y2=0
cc_247 N_B_c_281_n N_VGND_c_502_n 0.0105573f $X=2.52 $Y=0.18 $X2=0 $Y2=0
cc_248 N_B_M1009_g N_A_504_119#_c_551_n 0.0104018f $X=2.445 $Y=0.915 $X2=0 $Y2=0
cc_249 B N_A_504_119#_c_551_n 0.0198686f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_250 N_B_c_286_n N_A_504_119#_c_551_n 0.00134053f $X=2.42 $Y=1.51 $X2=0 $Y2=0
cc_251 N_B_c_280_n N_A_504_119#_c_552_n 0.0160463f $X=3.75 $Y=0.18 $X2=0 $Y2=0
cc_252 N_B_M1011_g N_A_504_119#_c_552_n 0.00390044f $X=3.825 $Y=0.915 $X2=0
+ $Y2=0
cc_253 N_B_M1009_g N_A_504_119#_c_553_n 0.00591191f $X=2.445 $Y=0.915 $X2=0
+ $Y2=0
cc_254 N_B_c_280_n N_A_504_119#_c_553_n 0.00778341f $X=3.75 $Y=0.18 $X2=0 $Y2=0
cc_255 N_B_c_281_n N_A_504_119#_c_553_n 2.14148e-19 $X=2.52 $Y=0.18 $X2=0 $Y2=0
cc_256 N_B_M1011_g N_A_504_119#_c_554_n 0.00289528f $X=3.825 $Y=0.915 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_356_n N_X_c_430_n 0.0691153f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_258 N_VPWR_c_357_n N_X_c_430_n 0.0525583f $X=1.18 $Y=2.35 $X2=0 $Y2=0
cc_259 N_VPWR_c_362_n N_X_c_430_n 0.0118568f $X=1.015 $Y=3.33 $X2=0 $Y2=0
cc_260 N_VPWR_c_354_n N_X_c_430_n 0.00973414f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_261 N_VPWR_M1012_d N_X_c_442_n 0.0037816f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_262 N_VPWR_c_357_n N_X_c_442_n 0.0154248f $X=1.18 $Y=2.35 $X2=0 $Y2=0
cc_263 N_VPWR_c_357_n N_X_c_431_n 0.0522442f $X=1.18 $Y=2.35 $X2=0 $Y2=0
cc_264 N_VPWR_c_358_n N_X_c_431_n 0.0430356f $X=2.1 $Y=2.455 $X2=0 $Y2=0
cc_265 N_VPWR_c_364_n N_X_c_431_n 0.0110241f $X=1.935 $Y=3.33 $X2=0 $Y2=0
cc_266 N_VPWR_c_354_n N_X_c_431_n 0.00909194f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_267 N_VPWR_c_356_n N_X_c_458_n 0.0131326f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_268 N_VPWR_c_356_n X 0.00179399f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_269 N_VPWR_c_356_n N_VGND_c_492_n 0.0100404f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_270 N_X_c_437_n N_VGND_M1004_d 0.00330483f $X=1.475 $Y=1.09 $X2=0 $Y2=0
cc_271 N_X_c_427_n N_VGND_c_492_n 0.0188983f $X=0.71 $Y=0.64 $X2=0 $Y2=0
cc_272 N_X_c_429_n N_VGND_c_492_n 0.0034415f $X=0.69 $Y=1.55 $X2=0 $Y2=0
cc_273 N_X_c_427_n N_VGND_c_493_n 0.0136308f $X=0.71 $Y=0.64 $X2=0 $Y2=0
cc_274 N_X_c_437_n N_VGND_c_493_n 0.0170777f $X=1.475 $Y=1.09 $X2=0 $Y2=0
cc_275 N_X_c_428_n N_VGND_c_493_n 0.014266f $X=1.64 $Y=0.64 $X2=0 $Y2=0
cc_276 N_X_c_437_n N_VGND_c_494_n 0.0101261f $X=1.475 $Y=1.09 $X2=0 $Y2=0
cc_277 N_X_c_428_n N_VGND_c_494_n 0.0290738f $X=1.64 $Y=0.64 $X2=0 $Y2=0
cc_278 N_X_c_427_n N_VGND_c_497_n 0.00727191f $X=0.71 $Y=0.64 $X2=0 $Y2=0
cc_279 N_X_c_428_n N_VGND_c_498_n 0.00734888f $X=1.64 $Y=0.64 $X2=0 $Y2=0
cc_280 N_X_c_427_n N_VGND_c_502_n 0.00841816f $X=0.71 $Y=0.64 $X2=0 $Y2=0
cc_281 N_X_c_428_n N_VGND_c_502_n 0.00845298f $X=1.64 $Y=0.64 $X2=0 $Y2=0
cc_282 N_VGND_c_494_n N_A_504_119#_c_551_n 0.0335983f $X=2.15 $Y=0.7 $X2=0 $Y2=0
cc_283 N_VGND_c_496_n N_A_504_119#_c_552_n 0.0126545f $X=4.04 $Y=0.74 $X2=0
+ $Y2=0
cc_284 N_VGND_c_499_n N_A_504_119#_c_552_n 0.0553269f $X=3.875 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_502_n N_A_504_119#_c_552_n 0.0286814f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_494_n N_A_504_119#_c_553_n 0.013618f $X=2.15 $Y=0.7 $X2=0 $Y2=0
cc_287 N_VGND_c_499_n N_A_504_119#_c_553_n 0.0224642f $X=3.875 $Y=0 $X2=0 $Y2=0
cc_288 N_VGND_c_502_n N_A_504_119#_c_553_n 0.0112854f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_289 N_VGND_c_496_n N_A_504_119#_c_554_n 0.0337444f $X=4.04 $Y=0.74 $X2=0
+ $Y2=0
