* NGSPICE file created from sky130_fd_sc_hs__a311o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 X a_154_392# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=1.947e+12p ps=1.641e+07u
M1001 VGND B1 a_154_392# VNB nlowvt w=640000u l=150000u
+  ad=1.23862e+12p pd=1.191e+07u as=5.376e+11p ps=5.52e+06u
M1002 VGND a_154_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1003 VPWR a_154_392# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_154_392# A1 a_1081_39# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=6.927e+11p ps=6.48e+06u
M1005 a_1081_39# A1 a_154_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_154_392# C1 a_69_392# VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=8.5e+11p ps=7.7e+06u
M1007 a_69_392# C1 a_154_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_154_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_888_105# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1010 a_1081_39# A2 a_888_105# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A3 a_888_105# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_334_392# B1 a_69_392# VPB pshort w=1e+06u l=150000u
+  ad=1.2e+12p pd=1.04e+07u as=0p ps=0u
M1013 a_334_392# A3 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND C1 a_154_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_154_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_334_392# A2 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A2 a_334_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_69_392# B1 a_334_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_888_105# A2 a_1081_39# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_154_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A3 a_334_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_334_392# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_154_392# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A1 a_334_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_154_392# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_154_392# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_154_392# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

