* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR RESET_B a_284_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X1 a_1429_308# a_1074_88# a_1827_144# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_2492_424# a_1827_144# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X3 VPWR a_854_74# a_1074_88# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 a_284_464# a_854_74# a_1272_131# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X5 a_324_81# D a_284_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_284_464# SCE a_538_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 VGND a_1272_131# a_1429_308# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_284_464# a_1074_88# a_1272_131# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 VPWR a_1272_131# a_1429_308# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 a_2087_410# a_1827_144# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 a_1827_144# a_1074_88# a_2073_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 VPWR a_2492_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 VPWR SCE a_206_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X14 a_1489_131# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 a_2492_424# a_1827_144# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X16 a_2265_74# a_1827_144# a_2087_410# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 VGND a_2492_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VPWR RESET_B a_1272_131# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X19 a_1272_131# a_854_74# a_1411_131# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 VGND RESET_B a_2265_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 VPWR CLK_N a_854_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X22 a_1429_308# a_854_74# a_1827_144# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 a_1827_144# a_854_74# a_2042_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X24 a_2042_508# a_2087_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X25 a_206_464# D a_284_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X26 a_471_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X27 a_1272_131# a_1074_88# a_1384_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X28 VPWR RESET_B a_2087_410# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X29 a_27_88# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X30 a_239_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 a_1411_131# a_1429_308# a_1489_131# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 a_239_81# a_27_88# a_324_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 a_538_81# SCD a_239_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 VGND a_854_74# a_1074_88# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 a_27_88# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 VGND CLK_N a_854_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 a_1384_508# a_1429_308# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X38 a_2073_74# a_2087_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 a_284_464# a_27_88# a_471_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
.ends
