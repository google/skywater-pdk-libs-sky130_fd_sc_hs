* File: sky130_fd_sc_hs__o311ai_4.spice
* Created: Thu Aug 27 21:02:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o311ai_4.pex.spice"
.subckt sky130_fd_sc_hs__o311ai_4  VNB VPB C1 B1 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1004 N_Y_M1004_d N_C1_M1004_g N_A_27_74#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.2109 PD=1.025 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1023 N_Y_M1004_d N_C1_M1023_g N_A_27_74#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1025 N_Y_M1025_d N_C1_M1025_g N_A_27_74#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1034 N_Y_M1025_d N_C1_M1034_g N_A_27_74#_M1034_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1002 N_A_459_74#_M1002_d N_B1_M1002_g N_A_27_74#_M1034_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1019 N_A_459_74#_M1002_d N_B1_M1019_g N_A_27_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1020 N_A_459_74#_M1020_d N_B1_M1020_g N_A_27_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1032 N_A_459_74#_M1020_d N_B1_M1032_g N_A_27_74#_M1032_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1073 AS=0.19515 PD=1.03 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75003.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A3_M1015_g N_A_459_74#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.19445 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75006 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A3_M1017_g N_A_459_74#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1773 AS=0.1036 PD=1.28 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75005.5 A=0.111 P=1.78 MULT=1
MM1029 N_VGND_M1017_d N_A3_M1029_g N_A_459_74#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1773 AS=0.1036 PD=1.28 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1035 N_VGND_M1035_d N_A3_M1035_g N_A_459_74#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1815 AS=0.1036 PD=1.29 PS=1.02 NRD=14.592 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1035_d N_A2_M1003_g N_A_459_74#_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1815 AS=0.1036 PD=1.29 PS=1.02 NRD=14.592 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_459_74#_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.7
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1005_d N_A2_M1021_g N_A_459_74#_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.13135 PD=1.06 PS=1.095 NRD=6.48 NRS=12.156 M=1 R=4.93333
+ SA=75003.1 SB=75003 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1030_d N_A2_M1030_g N_A_459_74#_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.13135 PD=1.02 PS=1.095 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1030_d N_A1_M1000_g N_A_459_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.1
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A1_M1001_g N_A_459_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.31265 AS=0.1036 PD=1.585 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.5
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1001_d N_A1_M1006_g N_A_459_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.31265 AS=0.10915 PD=1.585 PS=1.035 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75005.5 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A1_M1018_g N_A_459_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.10915 PD=2.05 PS=1.035 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_C1_M1008_g N_Y_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.294 PD=2.83 PS=1.645 NRD=1.7533 NRS=32.5247 M=1 R=7.46667
+ SA=75000.2 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1026 N_VPWR_M1026_d N_C1_M1026_g N_Y_M1008_s VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.294 PD=1.47 PS=1.645 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75000.9
+ SB=75002.6 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g N_VPWR_M1026_d VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75001.4
+ SB=75002.1 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1007_d N_B1_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=1.8984 PD=1.42 PS=5.63 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.8
+ SB=75001.6 A=0.168 P=2.54 MULT=1
MM1011 N_A_841_368#_M1011_d N_A3_M1011_g N_Y_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.2 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1022 N_A_841_368#_M1022_d N_A3_M1022_g N_Y_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2072 AS=0.196 PD=1.49 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.3 A=0.168 P=2.54 MULT=1
MM1027 N_A_841_368#_M1022_d N_A3_M1027_g N_Y_M1027_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2072 AS=0.2688 PD=1.49 PS=1.6 NRD=5.2599 NRS=7.0329 M=1 R=7.46667
+ SA=75001.2 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1028 N_A_841_368#_M1028_d N_A3_M1028_g N_Y_M1027_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2688 PD=1.42 PS=1.6 NRD=1.7533 NRS=28.1316 M=1 R=7.46667
+ SA=75001.9 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1010 N_A_1350_368#_M1010_d N_A2_M1010_g N_A_841_368#_M1028_d VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.3 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1012 N_A_1350_368#_M1010_d N_A2_M1012_g N_A_841_368#_M1012_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.224 PD=1.47 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.8 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1013 N_A_1350_368#_M1013_d N_A2_M1013_g N_A_841_368#_M1012_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1016 N_A_1350_368#_M1013_d N_A2_M1016_g N_A_841_368#_M1016_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.8 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1014 N_A_1350_368#_M1014_d N_A1_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1024 N_A_1350_368#_M1014_d N_A1_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1031 N_A_1350_368#_M1031_d N_A1_M1031_g N_VPWR_M1024_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1033 N_A_1350_368#_M1031_d N_A1_M1033_g N_VPWR_M1033_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX36_noxref VNB VPB NWDIODE A=21.2412 P=26.56
*
.include "sky130_fd_sc_hs__o311ai_4.pxi.spice"
*
.ends
*
*
