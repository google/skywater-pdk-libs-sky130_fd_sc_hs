* File: sky130_fd_sc_hs__a21boi_1.pex.spice
* Created: Thu Aug 27 20:24:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A21BOI_1%B1_N 1 2 3 5 6 8 10 11 12 13 19 20
r49 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.285
+ $Y=1.44 $X2=0.285 $Y2=1.44
r50 22 24 22.2462 $w=3.9e-07 $l=1.8e-07 $layer=POLY_cond $X=0.352 $Y=1.26
+ $X2=0.352 $Y2=1.44
r51 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.285
+ $Y=0.42 $X2=0.285 $Y2=0.42
r52 17 22 8.93446 $w=4.35e-07 $l=8.21584e-08 $layer=POLY_cond $X=0.337 $Y=1.185
+ $X2=0.352 $Y2=1.26
r53 17 19 97.8064 $w=4.35e-07 $l=7.65e-07 $layer=POLY_cond $X=0.337 $Y=1.185
+ $X2=0.337 $Y2=0.42
r54 13 25 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.285 $Y=1.295
+ $X2=0.285 $Y2=1.44
r55 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.285 $Y=0.925
+ $X2=0.285 $Y2=1.295
r56 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.285 $Y=0.555
+ $X2=0.285 $Y2=0.925
r57 11 20 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.285 $Y=0.555
+ $X2=0.285 $Y2=0.42
r58 8 10 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1 $Y=1.185 $X2=1
+ $Y2=0.835
r59 7 22 25.2441 $w=1.5e-07 $l=2.03e-07 $layer=POLY_cond $X=0.555 $Y=1.26
+ $X2=0.352 $Y2=1.26
r60 6 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=1.26
+ $X2=1 $Y2=1.185
r61 6 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.925 $Y=1.26
+ $X2=0.555 $Y2=1.26
r62 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=2.045
+ $X2=0.495 $Y2=2.54
r63 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=1.955 $X2=0.495
+ $Y2=2.045
r64 1 24 45.6156 $w=3.9e-07 $l=3.18575e-07 $layer=POLY_cond $X=0.495 $Y=1.695
+ $X2=0.352 $Y2=1.44
r65 1 2 101.065 $w=1.8e-07 $l=2.6e-07 $layer=POLY_cond $X=0.495 $Y=1.695
+ $X2=0.495 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_1%A_29_424# 1 2 7 9 10 12 15 17 18 21 24 26
+ 29 32 33
r69 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.385 $X2=1.45 $Y2=1.385
r70 27 33 0.588983 $w=3.3e-07 $l=1.03e-07 $layer=LI1_cond $X=0.95 $Y=1.385
+ $X2=0.847 $Y2=1.385
r71 27 29 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.95 $Y=1.385 $X2=1.45
+ $Y2=1.385
r72 25 33 8.03064 $w=1.87e-07 $l=1.73292e-07 $layer=LI1_cond $X=0.83 $Y=1.55
+ $X2=0.847 $Y2=1.385
r73 25 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.83 $Y=1.55
+ $X2=0.83 $Y2=1.775
r74 24 33 8.03064 $w=1.87e-07 $l=1.65e-07 $layer=LI1_cond $X=0.847 $Y=1.22
+ $X2=0.847 $Y2=1.385
r75 24 32 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=0.847 $Y=1.22
+ $X2=0.847 $Y2=1.05
r76 19 32 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=0.885
+ $X2=0.785 $Y2=1.05
r77 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.785 $Y=0.885
+ $X2=0.785 $Y2=0.795
r78 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.745 $Y=1.86
+ $X2=0.83 $Y2=1.775
r79 17 18 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.745 $Y=1.86
+ $X2=0.435 $Y2=1.86
r80 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.27 $Y=1.945
+ $X2=0.435 $Y2=1.86
r81 13 15 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.27 $Y=1.945
+ $X2=0.27 $Y2=2.265
r82 10 30 38.8445 $w=3.55e-07 $l=2.31571e-07 $layer=POLY_cond $X=1.68 $Y=1.22
+ $X2=1.52 $Y2=1.385
r83 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.68 $Y=1.22 $X2=1.68
+ $Y2=0.74
r84 7 30 68.0361 $w=3.55e-07 $l=4.46654e-07 $layer=POLY_cond $X=1.665 $Y=1.765
+ $X2=1.52 $Y2=1.385
r85 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.665 $Y=1.765
+ $X2=1.665 $Y2=2.4
r86 2 15 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=2.12 $X2=0.27 $Y2=2.265
r87 1 21 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.56 $X2=0.785 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_1%A1 3 5 7 8 12
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r35 8 12 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=1.515
r36 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.115 $Y=1.765
+ $X2=2.13 $Y2=1.515
r37 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.115 $Y=1.765
+ $X2=2.115 $Y2=2.4
r38 1 11 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.11 $Y=1.35
+ $X2=2.13 $Y2=1.515
r39 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.11 $Y=1.35 $X2=2.11
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_1%A2 1 3 4 6 7 8
r25 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.385 $X2=2.67 $Y2=1.385
r26 8 13 14.0162 $w=3.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.67 $Y2=1.365
r27 7 13 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.365 $X2=2.67
+ $Y2=1.365
r28 4 12 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.595 $Y=1.765
+ $X2=2.67 $Y2=1.385
r29 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.595 $Y=1.765
+ $X2=2.595 $Y2=2.4
r30 1 12 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.58 $Y=1.22
+ $X2=2.67 $Y2=1.385
r31 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.58 $Y=1.22 $X2=2.58
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
r36 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r42 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 25 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.76 $Y2=3.33
r44 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 20 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.76 $Y2=3.33
r48 20 22 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 16 30 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.19 $Y=3.33 $X2=2.16
+ $Y2=3.33
r52 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=3.33
+ $X2=2.355 $Y2=3.33
r53 15 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.52 $Y=3.33 $X2=3.12
+ $Y2=3.33
r54 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.52 $Y=3.33
+ $X2=2.355 $Y2=3.33
r55 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=3.245
+ $X2=2.355 $Y2=3.33
r56 11 13 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.355 $Y=3.245
+ $X2=2.355 $Y2=2.485
r57 7 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r58 7 9 44.4843 $w=2.48e-07 $l=9.65e-07 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=2.28
r59 2 13 300 $w=1.7e-07 $l=7.22807e-07 $layer=licon1_PDIFF $count=2 $X=2.19
+ $Y=1.84 $X2=2.355 $Y2=2.485
r60 1 9 300 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=2.12 $X2=0.72 $Y2=2.28
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_1%Y 1 2 7 10 13 16 17 18 19 23
r48 31 33 6.29226 $w=3.49e-07 $l=1.8e-07 $layer=LI1_cond $X=1.305 $Y=1.805
+ $X2=1.305 $Y2=1.985
r49 19 29 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=1.305 $Y=2.775
+ $X2=1.305 $Y2=2.815
r50 18 19 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.305 $Y=2.405
+ $X2=1.305 $Y2=2.775
r51 18 23 6.94085 $w=4.38e-07 $l=2.65e-07 $layer=LI1_cond $X=1.305 $Y=2.405
+ $X2=1.305 $Y2=2.14
r52 17 23 3.4677 $w=4.4e-07 $l=1.05e-07 $layer=LI1_cond $X=1.305 $Y=2.035
+ $X2=1.305 $Y2=2.14
r53 17 33 1.74785 $w=3.49e-07 $l=5e-08 $layer=LI1_cond $X=1.305 $Y=2.035
+ $X2=1.305 $Y2=1.985
r54 15 16 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.882 $Y=1.01
+ $X2=1.882 $Y2=1.18
r55 13 15 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.935 $Y=0.515
+ $X2=1.935 $Y2=1.01
r56 10 16 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.79 $Y=1.72
+ $X2=1.79 $Y2=1.18
r57 8 31 4.95691 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.525 $Y=1.805
+ $X2=1.305 $Y2=1.805
r58 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=1.805
+ $X2=1.79 $Y2=1.72
r59 7 8 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.705 $Y=1.805
+ $X2=1.525 $Y2=1.805
r60 2 33 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.44 $Y2=1.985
r61 2 29 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.44 $Y2=2.815
r62 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.755
+ $Y=0.37 $X2=1.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_1%A_348_368# 1 2 9 13 16 18
r25 20 21 3.12451 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=2.145
+ $X2=2.82 $Y2=2.23
r26 18 20 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.82 $Y=1.985
+ $X2=2.82 $Y2=2.145
r27 13 21 6.6412 $w=2.93e-07 $l=1.7e-07 $layer=LI1_cond $X=2.837 $Y=2.4
+ $X2=2.837 $Y2=2.23
r28 10 16 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.02 $Y=2.145
+ $X2=1.872 $Y2=2.145
r29 9 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=2.145
+ $X2=2.82 $Y2=2.145
r30 9 10 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.655 $Y=2.145
+ $X2=2.02 $Y2=2.145
r31 2 18 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.67
+ $Y=1.84 $X2=2.82 $Y2=1.985
r32 2 13 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=2.67
+ $Y=1.84 $X2=2.82 $Y2=2.4
r33 1 16 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.74
+ $Y=1.84 $X2=1.89 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_1%VGND 1 2 8 11 15 17 22 29 30 33 36
r39 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r42 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=2.795
+ $Y2=0
r44 27 29 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=3.12
+ $Y2=0
r45 23 33 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.375
+ $Y2=0
r46 23 25 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.68
+ $Y2=0
r47 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.795
+ $Y2=0
r48 22 25 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=1.68
+ $Y2=0
r49 20 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r50 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 17 33 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=1.375
+ $Y2=0
r52 17 19 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=0.24
+ $Y2=0
r53 15 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r54 15 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r55 15 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0
r57 9 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0.515
r58 8 14 2.62105 $w=5.1e-07 $l=9e-08 $layer=LI1_cond $X=1.375 $Y=0.505 $X2=1.375
+ $Y2=0.595
r59 7 33 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0
r60 7 8 9.85006 $w=5.08e-07 $l=4.2e-07 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0.505
r61 2 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.655
+ $Y=0.37 $X2=2.795 $Y2=0.515
r62 1 14 91 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.56 $X2=1.465 $Y2=0.595
.ends

