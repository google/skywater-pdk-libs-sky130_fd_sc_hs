* File: sky130_fd_sc_hs__and4b_4.pxi.spice
* Created: Tue Sep  1 19:56:13 2020
* 
x_PM_SKY130_FD_SC_HS__AND4B_4%A_N N_A_N_c_137_n N_A_N_M1012_g N_A_N_c_138_n
+ N_A_N_M1013_g A_N PM_SKY130_FD_SC_HS__AND4B_4%A_N
x_PM_SKY130_FD_SC_HS__AND4B_4%A_199_294# N_A_199_294#_M1014_s
+ N_A_199_294#_M1002_d N_A_199_294#_M1010_s N_A_199_294#_M1015_d
+ N_A_199_294#_M1021_s N_A_199_294#_c_169_n N_A_199_294#_M1001_g
+ N_A_199_294#_M1006_g N_A_199_294#_c_171_n N_A_199_294#_M1011_g
+ N_A_199_294#_c_180_n N_A_199_294#_M1007_g N_A_199_294#_c_181_n
+ N_A_199_294#_M1009_g N_A_199_294#_M1020_g N_A_199_294#_c_182_n
+ N_A_199_294#_M1023_g N_A_199_294#_M1024_g N_A_199_294#_c_175_n
+ N_A_199_294#_c_183_n N_A_199_294#_c_184_n N_A_199_294#_c_232_p
+ N_A_199_294#_c_176_n N_A_199_294#_c_177_n N_A_199_294#_c_217_p
+ N_A_199_294#_c_186_n N_A_199_294#_c_195_p N_A_199_294#_c_187_n
+ N_A_199_294#_c_178_n PM_SKY130_FD_SC_HS__AND4B_4%A_199_294#
x_PM_SKY130_FD_SC_HS__AND4B_4%D N_D_c_329_n N_D_M1005_g N_D_c_323_n N_D_c_331_n
+ N_D_M1010_g N_D_c_324_n N_D_M1008_g N_D_c_325_n N_D_M1018_g N_D_c_326_n D D D
+ N_D_c_328_n PM_SKY130_FD_SC_HS__AND4B_4%D
x_PM_SKY130_FD_SC_HS__AND4B_4%C N_C_c_383_n N_C_M1002_g N_C_c_384_n N_C_c_385_n
+ N_C_c_386_n N_C_M1000_g N_C_c_388_n N_C_c_395_n N_C_M1003_g N_C_M1016_g
+ N_C_c_390_n N_C_c_391_n N_C_c_392_n C N_C_c_393_n
+ PM_SKY130_FD_SC_HS__AND4B_4%C
x_PM_SKY130_FD_SC_HS__AND4B_4%A_27_368# N_A_27_368#_M1013_s N_A_27_368#_M1012_s
+ N_A_27_368#_M1014_g N_A_27_368#_c_474_n N_A_27_368#_M1019_g
+ N_A_27_368#_M1022_g N_A_27_368#_c_475_n N_A_27_368#_M1021_g
+ N_A_27_368#_c_466_n N_A_27_368#_c_476_n N_A_27_368#_c_485_n
+ N_A_27_368#_c_467_n N_A_27_368#_c_468_n N_A_27_368#_c_513_n
+ N_A_27_368#_c_469_n N_A_27_368#_c_470_n N_A_27_368#_c_478_n
+ N_A_27_368#_c_471_n N_A_27_368#_c_480_n N_A_27_368#_c_472_n
+ N_A_27_368#_c_473_n PM_SKY130_FD_SC_HS__AND4B_4%A_27_368#
x_PM_SKY130_FD_SC_HS__AND4B_4%B N_B_c_597_n N_B_c_598_n N_B_c_606_n N_B_M1015_g
+ N_B_M1004_g N_B_c_600_n N_B_c_601_n N_B_c_602_n N_B_M1025_g N_B_M1017_g B
+ PM_SKY130_FD_SC_HS__AND4B_4%B
x_PM_SKY130_FD_SC_HS__AND4B_4%VPWR N_VPWR_M1012_d N_VPWR_M1007_s N_VPWR_M1023_s
+ N_VPWR_M1005_d N_VPWR_M1003_s N_VPWR_M1019_d N_VPWR_M1025_s N_VPWR_c_664_n
+ N_VPWR_c_665_n N_VPWR_c_666_n N_VPWR_c_667_n N_VPWR_c_668_n N_VPWR_c_669_n
+ N_VPWR_c_670_n N_VPWR_c_671_n N_VPWR_c_672_n N_VPWR_c_673_n N_VPWR_c_674_n
+ N_VPWR_c_675_n N_VPWR_c_676_n VPWR N_VPWR_c_677_n N_VPWR_c_678_n
+ N_VPWR_c_679_n N_VPWR_c_680_n N_VPWR_c_681_n N_VPWR_c_682_n N_VPWR_c_663_n
+ PM_SKY130_FD_SC_HS__AND4B_4%VPWR
x_PM_SKY130_FD_SC_HS__AND4B_4%X N_X_M1006_s N_X_M1020_s N_X_M1001_d N_X_M1009_d
+ N_X_c_762_n N_X_c_757_n N_X_c_758_n X X X X X N_X_c_761_n X N_X_c_769_n
+ PM_SKY130_FD_SC_HS__AND4B_4%X
x_PM_SKY130_FD_SC_HS__AND4B_4%VGND N_VGND_M1013_d N_VGND_M1011_d N_VGND_M1024_d
+ N_VGND_M1008_d N_VGND_c_818_n N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n
+ N_VGND_c_822_n N_VGND_c_823_n N_VGND_c_824_n VGND N_VGND_c_825_n
+ N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n
+ N_VGND_c_831_n PM_SKY130_FD_SC_HS__AND4B_4%VGND
x_PM_SKY130_FD_SC_HS__AND4B_4%A_664_125# N_A_664_125#_M1000_d
+ N_A_664_125#_M1016_d N_A_664_125#_M1017_d N_A_664_125#_c_901_n
+ N_A_664_125#_c_902_n N_A_664_125#_c_903_n N_A_664_125#_c_904_n
+ N_A_664_125#_c_905_n N_A_664_125#_c_906_n N_A_664_125#_c_907_n
+ PM_SKY130_FD_SC_HS__AND4B_4%A_664_125#
x_PM_SKY130_FD_SC_HS__AND4B_4%A_751_125# N_A_751_125#_M1000_s
+ N_A_751_125#_M1018_s N_A_751_125#_c_961_n N_A_751_125#_c_963_n
+ N_A_751_125#_c_960_n PM_SKY130_FD_SC_HS__AND4B_4%A_751_125#
x_PM_SKY130_FD_SC_HS__AND4B_4%A_1136_125# N_A_1136_125#_M1004_s
+ N_A_1136_125#_M1022_d N_A_1136_125#_c_984_n N_A_1136_125#_c_985_n
+ N_A_1136_125#_c_986_n PM_SKY130_FD_SC_HS__AND4B_4%A_1136_125#
cc_1 VNB N_A_N_c_137_n 0.0449743f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_N_c_138_n 0.0208794f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.22
cc_3 VNB A_N 0.00916222f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_199_294#_c_169_n 0.0164758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_199_294#_M1006_g 0.0226641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_199_294#_c_171_n 0.00926078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_199_294#_M1011_g 0.0241832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_199_294#_M1020_g 0.0242295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_199_294#_M1024_g 0.0242307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_199_294#_c_175_n 0.00444332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_199_294#_c_176_n 0.00296626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_199_294#_c_177_n 0.00360386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_199_294#_c_178_n 0.0809608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_c_323_n 0.00884036f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.22
cc_15 VNB N_D_c_324_n 0.0148233f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.385
cc_16 VNB N_D_c_325_n 0.0142612f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.37
cc_17 VNB N_D_c_326_n 0.0050101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB D 0.010589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_D_c_328_n 0.0488578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_c_383_n 0.035618f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_21 VNB N_C_c_384_n 0.0655029f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.79
cc_22 VNB N_C_c_385_n 0.0223825f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.79
cc_23 VNB N_C_c_386_n 0.0124252f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_24 VNB N_C_M1000_g 0.0328565f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_25 VNB N_C_c_388_n 0.103403f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.37
cc_26 VNB N_C_M1016_g 0.0253364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C_c_390_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C_c_391_n 0.00839426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_C_c_392_n 0.0106507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_c_393_n 0.00341194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_368#_M1014_g 0.0185365f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.385
cc_32 VNB N_A_27_368#_M1022_g 0.0217497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_368#_c_466_n 0.02003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_368#_c_467_n 0.00244208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_368#_c_468_n 0.0182741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_368#_c_469_n 0.0170197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_368#_c_470_n 0.00646723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_368#_c_471_n 0.0297886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_368#_c_472_n 0.00142009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_368#_c_473_n 0.0213361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_B_c_597_n 0.00666875f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_42 VNB N_B_c_598_n 0.00994453f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_43 VNB N_B_M1004_g 0.0292859f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.385
cc_44 VNB N_B_c_600_n 0.104114f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_45 VNB N_B_c_601_n 0.00962308f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_46 VNB N_B_c_602_n 0.0187863f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.37
cc_47 VNB N_B_M1017_g 0.0363835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB B 0.00124747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VPWR_c_663_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_X_c_757_n 0.00596934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_X_c_758_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB X 0.00172508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB X 0.00280128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_X_c_761_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_818_n 0.0106049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_819_n 0.02097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_820_n 0.00987337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_821_n 0.0247003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_822_n 0.0102202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_823_n 0.0199677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_824_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_825_n 0.018718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_826_n 0.0356343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_827_n 0.0762007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_828_n 0.402809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_829_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_830_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_831_n 0.0043699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_664_125#_c_901_n 0.00708785f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.37
cc_70 VNB N_A_664_125#_c_902_n 0.0128721f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.37
cc_71 VNB N_A_664_125#_c_903_n 0.00493612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_664_125#_c_904_n 0.00385728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_664_125#_c_905_n 0.0382876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_664_125#_c_906_n 0.00335039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_664_125#_c_907_n 0.0213365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_751_125#_c_960_n 0.00273786f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.37
cc_77 VNB N_A_1136_125#_c_984_n 0.00255783f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_78 VNB N_A_1136_125#_c_985_n 0.00157665f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.385
cc_79 VNB N_A_1136_125#_c_986_n 0.00237075f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.37
cc_80 VPB N_A_N_c_137_n 0.0286753f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_81 VPB N_A_199_294#_c_169_n 0.0237478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_199_294#_c_180_n 0.015107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_199_294#_c_181_n 0.0159419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_199_294#_c_182_n 0.0162763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_199_294#_c_183_n 0.00139365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_199_294#_c_184_n 0.00602576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_199_294#_c_177_n 0.00297186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_199_294#_c_186_n 0.00346945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_199_294#_c_187_n 0.00872169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_199_294#_c_178_n 0.020194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_D_c_329_n 0.0166099f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_92 VPB N_D_c_323_n 0.0131155f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.22
cc_93 VPB N_D_c_331_n 0.0215772f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.79
cc_94 VPB N_D_c_326_n 0.0110139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB D 0.00260186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_D_c_328_n 0.0350186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_C_c_383_n 0.0344947f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_98 VPB N_C_c_395_n 0.0335317f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.37
cc_99 VPB N_C_c_391_n 0.00370107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_C_c_393_n 0.00311035f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_368#_c_474_n 0.0149714f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.385
cc_102 VPB N_A_27_368#_c_475_n 0.0154105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_368#_c_476_n 0.0153183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_368#_c_469_n 0.0146491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_27_368#_c_478_n 0.01385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_27_368#_c_471_n 0.00777552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_368#_c_480_n 0.0222378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_368#_c_472_n 0.00172979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_368#_c_473_n 0.0302056f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_B_c_598_n 0.00768018f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_111 VPB N_B_c_606_n 0.0212976f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_112 VPB N_B_c_602_n 0.0398633f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.37
cc_113 VPB B 9.29746e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_664_n 0.0109061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_665_n 0.00329267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_666_n 0.0212593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_667_n 0.00683921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_668_n 0.00667347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_669_n 0.00329222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_670_n 0.00261656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_671_n 0.0234846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_672_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_673_n 0.0355792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_674_n 0.0063829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_675_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_676_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_677_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_678_n 0.017758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_679_n 0.0276255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_680_n 0.00656601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_681_n 0.00643005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_682_n 0.0389631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_663_n 0.0827444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_X_c_762_n 0.00597179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB X 0.0015499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 N_A_N_c_137_n N_A_199_294#_c_169_n 0.0373909f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_137 A_N N_A_199_294#_c_169_n 5.51989e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A_N_c_137_n N_A_199_294#_M1006_g 0.0120427f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_N_c_138_n N_A_199_294#_M1006_g 0.0135044f $X=0.535 $Y=1.22 $X2=0
+ $Y2=0
cc_140 A_N N_A_199_294#_M1006_g 0.00213771f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A_N_c_138_n N_A_27_368#_c_466_n 0.00351224f $X=0.535 $Y=1.22 $X2=0
+ $Y2=0
cc_142 N_A_N_c_137_n N_A_27_368#_c_476_n 0.00759254f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_N_c_137_n N_A_27_368#_c_485_n 0.0141676f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_A_N_c_137_n N_A_27_368#_c_478_n 0.004814f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_145 A_N N_A_27_368#_c_478_n 0.00107599f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A_N_c_137_n N_A_27_368#_c_471_n 0.0152937f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_N_c_138_n N_A_27_368#_c_471_n 0.00417267f $X=0.535 $Y=1.22 $X2=0
+ $Y2=0
cc_148 A_N N_A_27_368#_c_471_n 0.0276149f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A_N_c_137_n N_A_27_368#_c_480_n 0.00607645f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_150 N_A_N_c_137_n N_VPWR_c_664_n 0.00446259f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_N_c_137_n N_VPWR_c_679_n 0.00481995f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_N_c_137_n N_VPWR_c_663_n 0.00508379f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_N_c_138_n X 4.11144e-19 $X=0.535 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A_N_c_137_n X 0.00167618f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_N_c_138_n X 2.30211e-19 $X=0.535 $Y=1.22 $X2=0 $Y2=0
cc_156 A_N X 0.0211453f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A_N_c_138_n N_X_c_761_n 2.11176e-19 $X=0.535 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A_N_c_137_n N_X_c_769_n 0.00135252f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_N_c_137_n N_VGND_c_818_n 8.95272e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A_N_c_138_n N_VGND_c_818_n 0.0135392f $X=0.535 $Y=1.22 $X2=0 $Y2=0
cc_161 A_N N_VGND_c_818_n 0.0189574f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_162 N_A_N_c_138_n N_VGND_c_825_n 0.00421418f $X=0.535 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A_N_c_138_n N_VGND_c_828_n 0.00432128f $X=0.535 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A_199_294#_c_186_n N_D_c_329_n 0.00136467f $X=3.515 $Y=2.085 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_199_294#_c_195_p N_D_c_329_n 0.0118815f $X=5.65 $Y=2.08 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A_199_294#_c_195_p N_D_c_323_n 0.00800297f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_167 N_A_199_294#_c_195_p N_D_c_331_n 0.0114222f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_168 N_A_199_294#_c_186_n N_D_c_326_n 4.55877e-19 $X=3.515 $Y=2.085 $X2=0
+ $Y2=0
cc_169 N_A_199_294#_c_195_p D 0.0842458f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_170 N_A_199_294#_c_195_p N_D_c_328_n 0.0141439f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_171 N_A_199_294#_c_182_n N_C_c_383_n 0.033124f $X=2.575 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A_199_294#_c_175_n N_C_c_383_n 0.00199938f $X=2.575 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_199_294#_c_183_n N_C_c_383_n 0.00360264f $X=2.66 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_199_294#_c_184_n N_C_c_383_n 0.0138403f $X=3.38 $Y=2.085 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_199_294#_c_178_n N_C_c_383_n 0.0191848f $X=2.575 $Y=1.542 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_199_294#_c_175_n N_C_c_384_n 7.00615e-19 $X=2.575 $Y=1.485 $X2=0
+ $Y2=0
cc_177 N_A_199_294#_c_178_n N_C_c_384_n 0.0116202f $X=2.575 $Y=1.542 $X2=0 $Y2=0
cc_178 N_A_199_294#_M1024_g N_C_c_386_n 0.0116202f $X=2.59 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_199_294#_c_195_p N_C_c_395_n 0.0114729f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_180 N_A_199_294#_c_175_n N_C_c_393_n 0.0253f $X=2.575 $Y=1.485 $X2=0 $Y2=0
cc_181 N_A_199_294#_c_183_n N_C_c_393_n 0.010144f $X=2.66 $Y=1.95 $X2=0 $Y2=0
cc_182 N_A_199_294#_c_184_n N_C_c_393_n 0.0262176f $X=3.38 $Y=2.085 $X2=0 $Y2=0
cc_183 N_A_199_294#_c_178_n N_C_c_393_n 6.22486e-19 $X=2.575 $Y=1.542 $X2=0
+ $Y2=0
cc_184 N_A_199_294#_c_176_n N_A_27_368#_M1014_g 0.0108741f $X=5.995 $Y=1.3 $X2=0
+ $Y2=0
cc_185 N_A_199_294#_c_177_n N_A_27_368#_M1014_g 0.00444636f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_186 N_A_199_294#_c_177_n N_A_27_368#_c_474_n 0.0019501f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_187 N_A_199_294#_c_217_p N_A_27_368#_c_474_n 0.00537234f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_188 N_A_199_294#_c_187_n N_A_27_368#_c_474_n 0.00558716f $X=6.08 $Y=2.08
+ $X2=0 $Y2=0
cc_189 N_A_199_294#_c_176_n N_A_27_368#_M1022_g 2.63345e-19 $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_190 N_A_199_294#_c_177_n N_A_27_368#_M1022_g 5.77979e-19 $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_191 N_A_199_294#_c_177_n N_A_27_368#_c_475_n 3.12965e-19 $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_192 N_A_199_294#_c_217_p N_A_27_368#_c_475_n 0.010767f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_193 N_A_199_294#_M1002_d N_A_27_368#_c_485_n 0.00549507f $X=3.2 $Y=1.96 $X2=0
+ $Y2=0
cc_194 N_A_199_294#_M1010_s N_A_27_368#_c_485_n 0.0262126f $X=4.185 $Y=1.96
+ $X2=0 $Y2=0
cc_195 N_A_199_294#_M1015_d N_A_27_368#_c_485_n 0.00549507f $X=5.665 $Y=1.96
+ $X2=0 $Y2=0
cc_196 N_A_199_294#_M1021_s N_A_27_368#_c_485_n 0.00549507f $X=6.565 $Y=1.96
+ $X2=0 $Y2=0
cc_197 N_A_199_294#_c_169_n N_A_27_368#_c_485_n 0.0146342f $X=1.085 $Y=1.765
+ $X2=0 $Y2=0
cc_198 N_A_199_294#_c_180_n N_A_27_368#_c_485_n 0.0119597f $X=1.535 $Y=1.765
+ $X2=0 $Y2=0
cc_199 N_A_199_294#_c_181_n N_A_27_368#_c_485_n 0.012516f $X=2.015 $Y=1.765
+ $X2=0 $Y2=0
cc_200 N_A_199_294#_c_182_n N_A_27_368#_c_485_n 0.0150655f $X=2.575 $Y=1.765
+ $X2=0 $Y2=0
cc_201 N_A_199_294#_c_184_n N_A_27_368#_c_485_n 0.240012f $X=3.38 $Y=2.085 $X2=0
+ $Y2=0
cc_202 N_A_199_294#_c_232_p N_A_27_368#_c_485_n 0.00871776f $X=2.745 $Y=2.085
+ $X2=0 $Y2=0
cc_203 N_A_199_294#_c_177_n N_A_27_368#_c_467_n 0.00543065f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_204 N_A_199_294#_c_217_p N_A_27_368#_c_468_n 0.00426251f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_205 N_A_199_294#_c_176_n N_A_27_368#_c_513_n 0.00867849f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_206 N_A_199_294#_c_217_p N_A_27_368#_c_469_n 0.00881186f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_207 N_A_199_294#_c_169_n N_A_27_368#_c_478_n 0.00197829f $X=1.085 $Y=1.765
+ $X2=0 $Y2=0
cc_208 N_A_199_294#_c_169_n N_A_27_368#_c_480_n 5.72061e-19 $X=1.085 $Y=1.765
+ $X2=0 $Y2=0
cc_209 N_A_199_294#_c_176_n N_A_27_368#_c_472_n 0.00681497f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_210 N_A_199_294#_c_177_n N_A_27_368#_c_472_n 0.0240318f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_211 N_A_199_294#_c_217_p N_A_27_368#_c_472_n 0.0278902f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_212 N_A_199_294#_c_176_n N_A_27_368#_c_473_n 0.00258046f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_213 N_A_199_294#_c_177_n N_A_27_368#_c_473_n 0.0132005f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_214 N_A_199_294#_c_217_p N_A_27_368#_c_473_n 0.00699607f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_215 N_A_199_294#_c_177_n N_B_c_606_n 0.00104603f $X=5.995 $Y=1.94 $X2=0 $Y2=0
cc_216 N_A_199_294#_c_195_p N_B_c_606_n 0.014386f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_217 N_A_199_294#_c_187_n N_B_c_606_n 0.00273592f $X=6.08 $Y=2.08 $X2=0 $Y2=0
cc_218 N_A_199_294#_c_176_n N_B_M1004_g 0.0011858f $X=5.995 $Y=1.3 $X2=0 $Y2=0
cc_219 N_A_199_294#_c_177_n N_B_M1004_g 0.0112606f $X=5.995 $Y=1.94 $X2=0 $Y2=0
cc_220 N_A_199_294#_c_217_p N_B_c_602_n 0.00472882f $X=6.715 $Y=2.135 $X2=0
+ $Y2=0
cc_221 N_A_199_294#_c_217_p B 0.00183728f $X=6.715 $Y=2.135 $X2=0 $Y2=0
cc_222 N_A_199_294#_c_183_n N_VPWR_M1023_s 0.00140032f $X=2.66 $Y=1.95 $X2=0
+ $Y2=0
cc_223 N_A_199_294#_c_184_n N_VPWR_M1023_s 0.010075f $X=3.38 $Y=2.085 $X2=0
+ $Y2=0
cc_224 N_A_199_294#_c_232_p N_VPWR_M1023_s 4.10458e-19 $X=2.745 $Y=2.085 $X2=0
+ $Y2=0
cc_225 N_A_199_294#_c_195_p N_VPWR_M1005_d 0.00722886f $X=5.65 $Y=2.08 $X2=0
+ $Y2=0
cc_226 N_A_199_294#_c_195_p N_VPWR_M1003_s 0.00662728f $X=5.65 $Y=2.08 $X2=0
+ $Y2=0
cc_227 N_A_199_294#_c_217_p N_VPWR_M1019_d 0.00401357f $X=6.715 $Y=2.135 $X2=0
+ $Y2=0
cc_228 N_A_199_294#_c_169_n N_VPWR_c_664_n 0.00941719f $X=1.085 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A_199_294#_c_180_n N_VPWR_c_664_n 0.00106388f $X=1.535 $Y=1.765 $X2=0
+ $Y2=0
cc_230 N_A_199_294#_c_169_n N_VPWR_c_665_n 0.00106413f $X=1.085 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_A_199_294#_c_180_n N_VPWR_c_665_n 0.00853363f $X=1.535 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_199_294#_c_181_n N_VPWR_c_665_n 0.00933219f $X=2.015 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A_199_294#_c_182_n N_VPWR_c_665_n 0.00163184f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A_199_294#_c_181_n N_VPWR_c_666_n 0.00413917f $X=2.015 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_A_199_294#_c_182_n N_VPWR_c_666_n 0.00413917f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A_199_294#_c_181_n N_VPWR_c_667_n 0.00163255f $X=2.015 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A_199_294#_c_182_n N_VPWR_c_667_n 0.00925933f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_199_294#_c_169_n N_VPWR_c_677_n 0.00413917f $X=1.085 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A_199_294#_c_180_n N_VPWR_c_677_n 0.00413917f $X=1.535 $Y=1.765 $X2=0
+ $Y2=0
cc_240 N_A_199_294#_c_169_n N_VPWR_c_663_n 0.00398641f $X=1.085 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A_199_294#_c_180_n N_VPWR_c_663_n 0.00398641f $X=1.535 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_A_199_294#_c_181_n N_VPWR_c_663_n 0.003996f $X=2.015 $Y=1.765 $X2=0
+ $Y2=0
cc_243 N_A_199_294#_c_182_n N_VPWR_c_663_n 0.003996f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A_199_294#_c_171_n N_X_c_762_n 8.03946e-19 $X=1.445 $Y=1.395 $X2=0
+ $Y2=0
cc_245 N_A_199_294#_c_180_n N_X_c_762_n 0.0158685f $X=1.535 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A_199_294#_c_181_n N_X_c_762_n 0.015525f $X=2.015 $Y=1.765 $X2=0 $Y2=0
cc_247 N_A_199_294#_c_182_n N_X_c_762_n 0.00355585f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A_199_294#_c_175_n N_X_c_762_n 0.0727822f $X=2.575 $Y=1.485 $X2=0 $Y2=0
cc_249 N_A_199_294#_c_183_n N_X_c_762_n 0.0101811f $X=2.66 $Y=1.95 $X2=0 $Y2=0
cc_250 N_A_199_294#_c_232_p N_X_c_762_n 0.0235115f $X=2.745 $Y=2.085 $X2=0 $Y2=0
cc_251 N_A_199_294#_c_178_n N_X_c_762_n 0.0167559f $X=2.575 $Y=1.542 $X2=0 $Y2=0
cc_252 N_A_199_294#_M1011_g N_X_c_757_n 0.0123455f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_199_294#_M1020_g N_X_c_757_n 0.0133553f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_199_294#_M1024_g N_X_c_757_n 0.00283169f $X=2.59 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_199_294#_c_175_n N_X_c_757_n 0.0811859f $X=2.575 $Y=1.485 $X2=0 $Y2=0
cc_256 N_A_199_294#_c_178_n N_X_c_757_n 0.00951805f $X=2.575 $Y=1.542 $X2=0
+ $Y2=0
cc_257 N_A_199_294#_M1011_g N_X_c_758_n 8.39752e-19 $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_199_294#_M1020_g N_X_c_758_n 0.010036f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_199_294#_M1024_g N_X_c_758_n 0.00768257f $X=2.59 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_199_294#_M1006_g X 0.00437707f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_199_294#_c_171_n X 0.00107372f $X=1.445 $Y=1.395 $X2=0 $Y2=0
cc_262 N_A_199_294#_M1011_g X 0.00153926f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_199_294#_c_169_n X 0.0132265f $X=1.085 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_199_294#_M1006_g X 0.004196f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_199_294#_c_171_n X 0.00662179f $X=1.445 $Y=1.395 $X2=0 $Y2=0
cc_266 N_A_199_294#_M1011_g X 0.00389182f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_199_294#_c_180_n X 0.00123283f $X=1.535 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A_199_294#_c_175_n X 0.0262135f $X=2.575 $Y=1.485 $X2=0 $Y2=0
cc_269 N_A_199_294#_c_178_n X 0.00402611f $X=2.575 $Y=1.542 $X2=0 $Y2=0
cc_270 N_A_199_294#_M1006_g N_X_c_761_n 0.010518f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_199_294#_M1011_g N_X_c_761_n 0.00998276f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A_199_294#_M1020_g N_X_c_761_n 8.33931e-19 $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A_199_294#_c_169_n N_X_c_769_n 0.0107157f $X=1.085 $Y=1.765 $X2=0 $Y2=0
cc_274 N_A_199_294#_M1006_g N_VGND_c_818_n 0.00974391f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_275 N_A_199_294#_M1006_g N_VGND_c_819_n 0.00371957f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_276 N_A_199_294#_M1011_g N_VGND_c_819_n 0.00434272f $X=1.52 $Y=0.74 $X2=0
+ $Y2=0
cc_277 N_A_199_294#_M1011_g N_VGND_c_820_n 0.0077868f $X=1.52 $Y=0.74 $X2=0
+ $Y2=0
cc_278 N_A_199_294#_M1020_g N_VGND_c_820_n 0.00772705f $X=2.16 $Y=0.74 $X2=0
+ $Y2=0
cc_279 N_A_199_294#_M1024_g N_VGND_c_821_n 0.00815524f $X=2.59 $Y=0.74 $X2=0
+ $Y2=0
cc_280 N_A_199_294#_c_175_n N_VGND_c_821_n 0.00294321f $X=2.575 $Y=1.485 $X2=0
+ $Y2=0
cc_281 N_A_199_294#_M1020_g N_VGND_c_823_n 0.00434272f $X=2.16 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A_199_294#_M1024_g N_VGND_c_823_n 0.00434272f $X=2.59 $Y=0.74 $X2=0
+ $Y2=0
cc_283 N_A_199_294#_M1006_g N_VGND_c_828_n 0.00624491f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_284 N_A_199_294#_M1011_g N_VGND_c_828_n 0.00822469f $X=1.52 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_199_294#_M1020_g N_VGND_c_828_n 0.00822693f $X=2.16 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_A_199_294#_M1024_g N_VGND_c_828_n 0.00821384f $X=2.59 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_199_294#_c_176_n N_A_664_125#_c_902_n 0.00159069f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_288 N_A_199_294#_c_195_p N_A_664_125#_c_902_n 0.0161891f $X=5.65 $Y=2.08
+ $X2=0 $Y2=0
cc_289 N_A_199_294#_c_186_n N_A_664_125#_c_903_n 0.00181215f $X=3.515 $Y=2.085
+ $X2=0 $Y2=0
cc_290 N_A_199_294#_c_195_p N_A_664_125#_c_903_n 0.00323763f $X=5.65 $Y=2.08
+ $X2=0 $Y2=0
cc_291 N_A_199_294#_M1014_s N_A_1136_125#_c_984_n 0.00176461f $X=6.11 $Y=0.625
+ $X2=0 $Y2=0
cc_292 N_A_199_294#_c_176_n N_A_1136_125#_c_984_n 0.0198997f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_293 N_D_c_329_n N_C_c_383_n 0.0360121f $X=3.575 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_294 N_D_c_326_n N_C_c_383_n 0.012499f $X=3.575 $Y=1.725 $X2=-0.19 $Y2=-0.245
cc_295 N_D_c_324_n N_C_M1000_g 0.0213925f $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_296 N_D_c_326_n N_C_M1000_g 0.00823494f $X=3.575 $Y=1.725 $X2=0 $Y2=0
cc_297 N_D_c_324_n N_C_c_388_n 0.00852785f $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_298 N_D_c_325_n N_C_c_388_n 0.00852641f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_299 D N_C_c_395_n 0.00478751f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_300 N_D_c_328_n N_C_c_395_n 0.00296558f $X=4.585 $Y=1.635 $X2=0 $Y2=0
cc_301 N_D_c_325_n N_C_M1016_g 0.0223678f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_302 D N_C_c_391_n 0.00914665f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_303 N_D_c_328_n N_C_c_391_n 0.0145538f $X=4.585 $Y=1.635 $X2=0 $Y2=0
cc_304 N_D_c_325_n N_C_c_392_n 0.00502045f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_305 D N_C_c_392_n 0.00179587f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_306 N_D_c_326_n N_C_c_393_n 0.00250476f $X=3.575 $Y=1.725 $X2=0 $Y2=0
cc_307 N_D_c_329_n N_A_27_368#_c_485_n 0.0122948f $X=3.575 $Y=1.885 $X2=0 $Y2=0
cc_308 N_D_c_331_n N_A_27_368#_c_485_n 0.0141558f $X=4.11 $Y=1.885 $X2=0 $Y2=0
cc_309 D N_B_c_597_n 0.00182248f $X=4.955 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_310 N_D_c_329_n N_VPWR_c_668_n 0.0100139f $X=3.575 $Y=1.885 $X2=0 $Y2=0
cc_311 N_D_c_331_n N_VPWR_c_668_n 0.0173454f $X=4.11 $Y=1.885 $X2=0 $Y2=0
cc_312 N_D_c_329_n N_VPWR_c_671_n 0.00461464f $X=3.575 $Y=1.885 $X2=0 $Y2=0
cc_313 N_D_c_331_n N_VPWR_c_673_n 0.00413917f $X=4.11 $Y=1.885 $X2=0 $Y2=0
cc_314 N_D_c_329_n N_VPWR_c_663_n 0.00447679f $X=3.575 $Y=1.885 $X2=0 $Y2=0
cc_315 N_D_c_331_n N_VPWR_c_663_n 0.00403443f $X=4.11 $Y=1.885 $X2=0 $Y2=0
cc_316 N_D_c_324_n N_VGND_c_822_n 0.00344336f $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_317 N_D_c_325_n N_VGND_c_822_n 0.00334294f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_318 N_D_c_324_n N_VGND_c_828_n 9.49986e-19 $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_319 N_D_c_325_n N_VGND_c_828_n 9.49986e-19 $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_320 N_D_c_324_n N_A_664_125#_c_901_n 8.29779e-19 $X=4.155 $Y=1.345 $X2=0
+ $Y2=0
cc_321 N_D_c_323_n N_A_664_125#_c_902_n 0.0045448f $X=4.02 $Y=1.725 $X2=0 $Y2=0
cc_322 N_D_c_324_n N_A_664_125#_c_902_n 0.0114991f $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_323 N_D_c_325_n N_A_664_125#_c_902_n 0.0112328f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_324 N_D_c_326_n N_A_664_125#_c_902_n 4.32292e-19 $X=3.575 $Y=1.725 $X2=0
+ $Y2=0
cc_325 D N_A_664_125#_c_902_n 0.0895722f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_326 N_D_c_328_n N_A_664_125#_c_902_n 0.00722393f $X=4.585 $Y=1.635 $X2=0
+ $Y2=0
cc_327 N_D_c_326_n N_A_664_125#_c_903_n 0.00329037f $X=3.575 $Y=1.725 $X2=0
+ $Y2=0
cc_328 N_D_c_324_n N_A_751_125#_c_961_n 0.00759913f $X=4.155 $Y=1.345 $X2=0
+ $Y2=0
cc_329 N_D_c_325_n N_A_751_125#_c_961_n 0.00813572f $X=4.745 $Y=1.345 $X2=0
+ $Y2=0
cc_330 N_D_c_324_n N_A_751_125#_c_963_n 0.00433778f $X=4.155 $Y=1.345 $X2=0
+ $Y2=0
cc_331 N_D_c_325_n N_A_751_125#_c_963_n 7.19935e-19 $X=4.745 $Y=1.345 $X2=0
+ $Y2=0
cc_332 N_D_c_324_n N_A_751_125#_c_960_n 8.5254e-19 $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_333 N_D_c_325_n N_A_751_125#_c_960_n 0.00545393f $X=4.745 $Y=1.345 $X2=0
+ $Y2=0
cc_334 N_C_c_383_n N_A_27_368#_c_485_n 0.0122949f $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_335 N_C_c_395_n N_A_27_368#_c_485_n 0.0137705f $X=5.12 $Y=1.885 $X2=0 $Y2=0
cc_336 N_C_c_392_n N_B_c_597_n 0.00513299f $X=5.155 $Y=1.49 $X2=-0.19 $Y2=-0.245
cc_337 N_C_c_391_n N_B_c_598_n 0.00893813f $X=5.12 $Y=1.735 $X2=0 $Y2=0
cc_338 N_C_c_395_n N_B_c_606_n 0.0437861f $X=5.12 $Y=1.885 $X2=0 $Y2=0
cc_339 N_C_M1016_g N_B_M1004_g 0.0138613f $X=5.175 $Y=0.945 $X2=0 $Y2=0
cc_340 N_C_c_388_n N_B_c_601_n 0.0138613f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_341 N_C_c_383_n N_VPWR_c_667_n 0.0101592f $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_342 N_C_c_395_n N_VPWR_c_669_n 0.0174676f $X=5.12 $Y=1.885 $X2=0 $Y2=0
cc_343 N_C_c_383_n N_VPWR_c_671_n 0.00461464f $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_344 N_C_c_395_n N_VPWR_c_673_n 0.00413917f $X=5.12 $Y=1.885 $X2=0 $Y2=0
cc_345 N_C_c_383_n N_VPWR_c_663_n 0.00447828f $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_346 N_C_c_395_n N_VPWR_c_663_n 0.00403443f $X=5.12 $Y=1.885 $X2=0 $Y2=0
cc_347 N_C_c_383_n N_VGND_c_821_n 9.4278e-19 $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_348 N_C_c_386_n N_VGND_c_821_n 0.0213937f $X=3.245 $Y=0.18 $X2=0 $Y2=0
cc_349 N_C_c_393_n N_VGND_c_821_n 0.008741f $X=3.08 $Y=1.515 $X2=0 $Y2=0
cc_350 N_C_M1000_g N_VGND_c_822_n 0.00634879f $X=3.68 $Y=0.945 $X2=0 $Y2=0
cc_351 N_C_c_388_n N_VGND_c_822_n 0.025075f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_352 N_C_M1016_g N_VGND_c_822_n 0.00659036f $X=5.175 $Y=0.945 $X2=0 $Y2=0
cc_353 N_C_c_386_n N_VGND_c_826_n 0.0372748f $X=3.245 $Y=0.18 $X2=0 $Y2=0
cc_354 N_C_c_388_n N_VGND_c_827_n 0.0196635f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_355 N_C_c_385_n N_VGND_c_828_n 0.0116023f $X=3.605 $Y=0.18 $X2=0 $Y2=0
cc_356 N_C_c_386_n N_VGND_c_828_n 0.011445f $X=3.245 $Y=0.18 $X2=0 $Y2=0
cc_357 N_C_c_388_n N_VGND_c_828_n 0.0386483f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_358 N_C_c_390_n N_VGND_c_828_n 0.00846253f $X=3.68 $Y=0.18 $X2=0 $Y2=0
cc_359 N_C_c_384_n N_A_664_125#_c_901_n 0.00523221f $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_360 N_C_c_385_n N_A_664_125#_c_901_n 0.00353352f $X=3.605 $Y=0.18 $X2=0 $Y2=0
cc_361 N_C_M1000_g N_A_664_125#_c_901_n 0.00930239f $X=3.68 $Y=0.945 $X2=0 $Y2=0
cc_362 N_C_M1000_g N_A_664_125#_c_902_n 0.0116916f $X=3.68 $Y=0.945 $X2=0 $Y2=0
cc_363 N_C_M1016_g N_A_664_125#_c_902_n 0.0136463f $X=5.175 $Y=0.945 $X2=0 $Y2=0
cc_364 N_C_c_392_n N_A_664_125#_c_902_n 0.00122885f $X=5.155 $Y=1.49 $X2=0 $Y2=0
cc_365 N_C_c_384_n N_A_664_125#_c_903_n 0.00485899f $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_366 N_C_M1000_g N_A_664_125#_c_903_n 0.00248638f $X=3.68 $Y=0.945 $X2=0 $Y2=0
cc_367 N_C_M1016_g N_A_664_125#_c_904_n 0.0044159f $X=5.175 $Y=0.945 $X2=0 $Y2=0
cc_368 N_C_M1016_g N_A_664_125#_c_906_n 0.00537518f $X=5.175 $Y=0.945 $X2=0
+ $Y2=0
cc_369 N_C_c_388_n N_A_751_125#_c_961_n 0.00200023f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_370 N_C_c_388_n N_A_751_125#_c_963_n 0.00413604f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_371 N_C_c_388_n N_A_751_125#_c_960_n 0.00367611f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_372 N_C_M1016_g N_A_751_125#_c_960_n 0.00469613f $X=5.175 $Y=0.945 $X2=0
+ $Y2=0
cc_373 N_A_27_368#_c_473_n N_B_c_597_n 0.0162934f $X=6.465 $Y=1.677 $X2=-0.19
+ $Y2=-0.245
cc_374 N_A_27_368#_c_473_n N_B_c_598_n 0.0116064f $X=6.465 $Y=1.677 $X2=0 $Y2=0
cc_375 N_A_27_368#_c_474_n N_B_c_606_n 0.0351028f $X=6.04 $Y=1.885 $X2=0 $Y2=0
cc_376 N_A_27_368#_c_485_n N_B_c_606_n 0.0117989f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_377 N_A_27_368#_M1014_g N_B_M1004_g 0.0162934f $X=6.035 $Y=0.945 $X2=0 $Y2=0
cc_378 N_A_27_368#_M1014_g N_B_c_600_n 0.00737859f $X=6.035 $Y=0.945 $X2=0 $Y2=0
cc_379 N_A_27_368#_M1022_g N_B_c_600_n 0.00737859f $X=6.465 $Y=0.945 $X2=0 $Y2=0
cc_380 N_A_27_368#_c_475_n N_B_c_602_n 0.0350555f $X=6.49 $Y=1.885 $X2=0 $Y2=0
cc_381 N_A_27_368#_c_485_n N_B_c_602_n 0.0181273f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_382 N_A_27_368#_c_468_n N_B_c_602_n 0.00488346f $X=7.35 $Y=1.215 $X2=0 $Y2=0
cc_383 N_A_27_368#_c_469_n N_B_c_602_n 0.0143843f $X=7.435 $Y=2.39 $X2=0 $Y2=0
cc_384 N_A_27_368#_c_472_n N_B_c_602_n 0.00117267f $X=6.59 $Y=1.635 $X2=0 $Y2=0
cc_385 N_A_27_368#_c_473_n N_B_c_602_n 0.0203498f $X=6.465 $Y=1.677 $X2=0 $Y2=0
cc_386 N_A_27_368#_M1022_g N_B_M1017_g 0.0182961f $X=6.465 $Y=0.945 $X2=0 $Y2=0
cc_387 N_A_27_368#_c_467_n N_B_M1017_g 7.10656e-19 $X=6.59 $Y=1.47 $X2=0 $Y2=0
cc_388 N_A_27_368#_c_468_n N_B_M1017_g 0.0170156f $X=7.35 $Y=1.215 $X2=0 $Y2=0
cc_389 N_A_27_368#_c_469_n N_B_M1017_g 0.0123314f $X=7.435 $Y=2.39 $X2=0 $Y2=0
cc_390 N_A_27_368#_c_485_n B 0.00721403f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_391 N_A_27_368#_c_468_n B 0.0246739f $X=7.35 $Y=1.215 $X2=0 $Y2=0
cc_392 N_A_27_368#_c_469_n B 0.0248009f $X=7.435 $Y=2.39 $X2=0 $Y2=0
cc_393 N_A_27_368#_c_472_n B 0.0281241f $X=6.59 $Y=1.635 $X2=0 $Y2=0
cc_394 N_A_27_368#_c_473_n B 9.04921e-19 $X=6.465 $Y=1.677 $X2=0 $Y2=0
cc_395 N_A_27_368#_c_485_n N_VPWR_M1012_d 0.0161195f $X=7.35 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_396 N_A_27_368#_c_485_n N_VPWR_M1007_s 0.00455255f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_397 N_A_27_368#_c_485_n N_VPWR_M1023_s 0.00649614f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_398 N_A_27_368#_c_485_n N_VPWR_M1005_d 0.00580876f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_399 N_A_27_368#_c_485_n N_VPWR_M1003_s 0.00434179f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_400 N_A_27_368#_c_485_n N_VPWR_M1019_d 0.00374591f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_401 N_A_27_368#_c_485_n N_VPWR_M1025_s 0.0234761f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_402 N_A_27_368#_c_469_n N_VPWR_M1025_s 0.0261656f $X=7.435 $Y=2.39 $X2=0
+ $Y2=0
cc_403 N_A_27_368#_c_485_n N_VPWR_c_664_n 0.0248792f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_404 N_A_27_368#_c_480_n N_VPWR_c_664_n 0.00891314f $X=0.265 $Y=2.475 $X2=0
+ $Y2=0
cc_405 N_A_27_368#_c_485_n N_VPWR_c_665_n 0.0190723f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_406 N_A_27_368#_c_485_n N_VPWR_c_667_n 0.0225065f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_407 N_A_27_368#_c_485_n N_VPWR_c_668_n 0.0213202f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_408 N_A_27_368#_c_474_n N_VPWR_c_669_n 0.0010643f $X=6.04 $Y=1.885 $X2=0
+ $Y2=0
cc_409 N_A_27_368#_c_485_n N_VPWR_c_669_n 0.0182814f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_410 N_A_27_368#_c_474_n N_VPWR_c_670_n 0.00840438f $X=6.04 $Y=1.885 $X2=0
+ $Y2=0
cc_411 N_A_27_368#_c_475_n N_VPWR_c_670_n 0.00839869f $X=6.49 $Y=1.885 $X2=0
+ $Y2=0
cc_412 N_A_27_368#_c_485_n N_VPWR_c_670_n 0.0166996f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_413 N_A_27_368#_c_474_n N_VPWR_c_675_n 0.00413917f $X=6.04 $Y=1.885 $X2=0
+ $Y2=0
cc_414 N_A_27_368#_c_475_n N_VPWR_c_678_n 0.00413917f $X=6.49 $Y=1.885 $X2=0
+ $Y2=0
cc_415 N_A_27_368#_c_480_n N_VPWR_c_679_n 0.0106977f $X=0.265 $Y=2.475 $X2=0
+ $Y2=0
cc_416 N_A_27_368#_c_475_n N_VPWR_c_682_n 0.00106308f $X=6.49 $Y=1.885 $X2=0
+ $Y2=0
cc_417 N_A_27_368#_c_485_n N_VPWR_c_682_n 0.0378332f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_418 N_A_27_368#_c_474_n N_VPWR_c_663_n 0.00398725f $X=6.04 $Y=1.885 $X2=0
+ $Y2=0
cc_419 N_A_27_368#_c_475_n N_VPWR_c_663_n 0.00398725f $X=6.49 $Y=1.885 $X2=0
+ $Y2=0
cc_420 N_A_27_368#_c_485_n N_VPWR_c_663_n 0.161342f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_421 N_A_27_368#_c_480_n N_VPWR_c_663_n 0.0122155f $X=0.265 $Y=2.475 $X2=0
+ $Y2=0
cc_422 N_A_27_368#_c_485_n N_X_M1001_d 0.00549253f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_423 N_A_27_368#_c_485_n N_X_M1009_d 0.0102548f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_424 N_A_27_368#_c_485_n N_X_c_762_n 0.0653239f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_425 N_A_27_368#_c_485_n N_X_c_769_n 0.0136442f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_426 N_A_27_368#_c_478_n N_X_c_769_n 0.0106116f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_427 N_A_27_368#_c_466_n N_VGND_c_818_n 0.0211853f $X=0.245 $Y=0.86 $X2=0
+ $Y2=0
cc_428 N_A_27_368#_c_466_n N_VGND_c_825_n 0.0100349f $X=0.245 $Y=0.86 $X2=0
+ $Y2=0
cc_429 N_A_27_368#_c_466_n N_VGND_c_828_n 0.0109771f $X=0.245 $Y=0.86 $X2=0
+ $Y2=0
cc_430 N_A_27_368#_c_468_n N_A_664_125#_M1017_d 0.00315946f $X=7.35 $Y=1.215
+ $X2=0 $Y2=0
cc_431 N_A_27_368#_M1014_g N_A_664_125#_c_905_n 0.00116683f $X=6.035 $Y=0.945
+ $X2=0 $Y2=0
cc_432 N_A_27_368#_M1022_g N_A_664_125#_c_905_n 0.00116683f $X=6.465 $Y=0.945
+ $X2=0 $Y2=0
cc_433 N_A_27_368#_M1022_g N_A_664_125#_c_907_n 5.83127e-19 $X=6.465 $Y=0.945
+ $X2=0 $Y2=0
cc_434 N_A_27_368#_c_468_n N_A_664_125#_c_907_n 0.023263f $X=7.35 $Y=1.215 $X2=0
+ $Y2=0
cc_435 N_A_27_368#_c_468_n N_A_1136_125#_M1022_d 0.00527828f $X=7.35 $Y=1.215
+ $X2=0 $Y2=0
cc_436 N_A_27_368#_c_513_n N_A_1136_125#_M1022_d 9.89161e-19 $X=6.675 $Y=1.215
+ $X2=0 $Y2=0
cc_437 N_A_27_368#_M1014_g N_A_1136_125#_c_984_n 0.00839754f $X=6.035 $Y=0.945
+ $X2=0 $Y2=0
cc_438 N_A_27_368#_M1022_g N_A_1136_125#_c_984_n 0.0128612f $X=6.465 $Y=0.945
+ $X2=0 $Y2=0
cc_439 N_A_27_368#_c_513_n N_A_1136_125#_c_984_n 0.00258843f $X=6.675 $Y=1.215
+ $X2=0 $Y2=0
cc_440 N_A_27_368#_M1022_g N_A_1136_125#_c_986_n 0.00532016f $X=6.465 $Y=0.945
+ $X2=0 $Y2=0
cc_441 N_A_27_368#_c_468_n N_A_1136_125#_c_986_n 0.0193536f $X=7.35 $Y=1.215
+ $X2=0 $Y2=0
cc_442 N_A_27_368#_c_513_n N_A_1136_125#_c_986_n 0.00360032f $X=6.675 $Y=1.215
+ $X2=0 $Y2=0
cc_443 N_B_c_606_n N_VPWR_c_669_n 0.00844933f $X=5.59 $Y=1.885 $X2=0 $Y2=0
cc_444 N_B_c_606_n N_VPWR_c_670_n 0.00106466f $X=5.59 $Y=1.885 $X2=0 $Y2=0
cc_445 N_B_c_602_n N_VPWR_c_670_n 0.00106425f $X=6.94 $Y=1.885 $X2=0 $Y2=0
cc_446 N_B_c_606_n N_VPWR_c_675_n 0.00413917f $X=5.59 $Y=1.885 $X2=0 $Y2=0
cc_447 N_B_c_602_n N_VPWR_c_678_n 0.00413917f $X=6.94 $Y=1.885 $X2=0 $Y2=0
cc_448 N_B_c_602_n N_VPWR_c_682_n 0.0151152f $X=6.94 $Y=1.885 $X2=0 $Y2=0
cc_449 N_B_c_606_n N_VPWR_c_663_n 0.00398725f $X=5.59 $Y=1.885 $X2=0 $Y2=0
cc_450 N_B_c_602_n N_VPWR_c_663_n 0.00397192f $X=6.94 $Y=1.885 $X2=0 $Y2=0
cc_451 N_B_c_601_n N_VGND_c_827_n 0.0351645f $X=5.68 $Y=0.18 $X2=0 $Y2=0
cc_452 N_B_c_600_n N_VGND_c_828_n 0.0374956f $X=7.04 $Y=0.18 $X2=0 $Y2=0
cc_453 N_B_c_601_n N_VGND_c_828_n 0.00460771f $X=5.68 $Y=0.18 $X2=0 $Y2=0
cc_454 N_B_M1004_g N_A_664_125#_c_902_n 4.46128e-19 $X=5.605 $Y=0.945 $X2=0
+ $Y2=0
cc_455 N_B_M1004_g N_A_664_125#_c_904_n 0.00424861f $X=5.605 $Y=0.945 $X2=0
+ $Y2=0
cc_456 N_B_M1004_g N_A_664_125#_c_905_n 0.0151367f $X=5.605 $Y=0.945 $X2=0 $Y2=0
cc_457 N_B_c_600_n N_A_664_125#_c_905_n 0.0230464f $X=7.04 $Y=0.18 $X2=0 $Y2=0
cc_458 N_B_M1017_g N_A_664_125#_c_905_n 0.0142293f $X=7.115 $Y=0.945 $X2=0 $Y2=0
cc_459 N_B_M1017_g N_A_664_125#_c_907_n 0.013896f $X=7.115 $Y=0.945 $X2=0 $Y2=0
cc_460 N_B_M1004_g N_A_1136_125#_c_985_n 0.00547385f $X=5.605 $Y=0.945 $X2=0
+ $Y2=0
cc_461 N_B_M1017_g N_A_1136_125#_c_986_n 0.00345017f $X=7.115 $Y=0.945 $X2=0
+ $Y2=0
cc_462 N_VPWR_M1007_s N_X_c_762_n 0.00236312f $X=1.61 $Y=1.84 $X2=0 $Y2=0
cc_463 N_X_c_757_n N_VGND_M1011_d 0.00624639f $X=2.21 $Y=1.065 $X2=0 $Y2=0
cc_464 X N_VGND_c_818_n 0.00329614f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_465 N_X_c_761_n N_VGND_c_818_n 0.0494597f $X=1.305 $Y=0.515 $X2=0 $Y2=0
cc_466 N_X_c_761_n N_VGND_c_819_n 0.0167819f $X=1.305 $Y=0.515 $X2=0 $Y2=0
cc_467 N_X_c_757_n N_VGND_c_820_n 0.0266856f $X=2.21 $Y=1.065 $X2=0 $Y2=0
cc_468 N_X_c_758_n N_VGND_c_820_n 0.0303828f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_469 N_X_c_761_n N_VGND_c_820_n 0.0319008f $X=1.305 $Y=0.515 $X2=0 $Y2=0
cc_470 N_X_c_757_n N_VGND_c_821_n 0.00711243f $X=2.21 $Y=1.065 $X2=0 $Y2=0
cc_471 N_X_c_758_n N_VGND_c_821_n 0.0243921f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_472 N_X_c_758_n N_VGND_c_823_n 0.0144922f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_473 N_X_c_758_n N_VGND_c_828_n 0.0118826f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_474 N_X_c_761_n N_VGND_c_828_n 0.0136487f $X=1.305 $Y=0.515 $X2=0 $Y2=0
cc_475 N_VGND_c_821_n N_A_664_125#_c_901_n 0.0324343f $X=2.875 $Y=0.515 $X2=0
+ $Y2=0
cc_476 N_VGND_c_822_n N_A_664_125#_c_901_n 4.21282e-19 $X=4.45 $Y=0.535 $X2=0
+ $Y2=0
cc_477 N_VGND_c_826_n N_A_664_125#_c_901_n 0.00697755f $X=4.285 $Y=0 $X2=0 $Y2=0
cc_478 N_VGND_c_828_n N_A_664_125#_c_901_n 0.00879953f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_479 N_VGND_M1008_d N_A_664_125#_c_902_n 0.00406725f $X=4.23 $Y=0.625 $X2=0
+ $Y2=0
cc_480 N_VGND_c_827_n N_A_664_125#_c_905_n 0.131618f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_481 N_VGND_c_828_n N_A_664_125#_c_905_n 0.0695304f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_482 N_VGND_c_827_n N_A_664_125#_c_906_n 0.0121867f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_828_n N_A_664_125#_c_906_n 0.00660921f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_484 N_VGND_M1008_d N_A_751_125#_c_961_n 0.00687044f $X=4.23 $Y=0.625 $X2=0
+ $Y2=0
cc_485 N_VGND_c_822_n N_A_751_125#_c_961_n 0.0260575f $X=4.45 $Y=0.535 $X2=0
+ $Y2=0
cc_486 N_VGND_c_828_n N_A_751_125#_c_961_n 0.0119525f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_c_826_n N_A_751_125#_c_963_n 0.00490296f $X=4.285 $Y=0 $X2=0 $Y2=0
cc_488 N_VGND_c_828_n N_A_751_125#_c_963_n 0.00747787f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_489 N_VGND_c_822_n N_A_751_125#_c_960_n 0.00113701f $X=4.45 $Y=0.535 $X2=0
+ $Y2=0
cc_490 N_VGND_c_827_n N_A_751_125#_c_960_n 0.00663395f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_491 N_VGND_c_828_n N_A_751_125#_c_960_n 0.00851925f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_492 N_A_664_125#_c_902_n N_A_751_125#_M1000_s 0.00224844f $X=5.305 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_493 N_A_664_125#_c_902_n N_A_751_125#_M1018_s 0.00176461f $X=5.305 $Y=1.215
+ $X2=0 $Y2=0
cc_494 N_A_664_125#_c_902_n N_A_751_125#_c_963_n 0.0584624f $X=5.305 $Y=1.215
+ $X2=0 $Y2=0
cc_495 N_A_664_125#_c_902_n N_A_751_125#_c_960_n 0.0162105f $X=5.305 $Y=1.215
+ $X2=0 $Y2=0
cc_496 N_A_664_125#_c_904_n N_A_751_125#_c_960_n 0.0134102f $X=5.39 $Y=0.77
+ $X2=0 $Y2=0
cc_497 N_A_664_125#_c_905_n N_A_1136_125#_c_984_n 0.0500146f $X=7.165 $Y=0.34
+ $X2=0 $Y2=0
cc_498 N_A_664_125#_c_904_n N_A_1136_125#_c_985_n 0.0135851f $X=5.39 $Y=0.77
+ $X2=0 $Y2=0
cc_499 N_A_664_125#_c_905_n N_A_1136_125#_c_985_n 0.0185025f $X=7.165 $Y=0.34
+ $X2=0 $Y2=0
cc_500 N_A_664_125#_c_905_n N_A_1136_125#_c_986_n 0.0245759f $X=7.165 $Y=0.34
+ $X2=0 $Y2=0
cc_501 N_A_664_125#_c_907_n N_A_1136_125#_c_986_n 0.0224808f $X=7.33 $Y=0.78
+ $X2=0 $Y2=0
