* NGSPICE file created from sky130_fd_sc_hs__and4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4_1 A B C D VGND VNB VPB VPWR X
M1000 VGND D a_335_74# VNB nlowvt w=640000u l=150000u
+  ad=2.554e+11p pd=2.2e+06u as=2.688e+11p ps=2.12e+06u
M1001 X a_96_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1002 VPWR B a_96_74# VPB pshort w=840000u l=150000u
+  ad=1.1998e+12p pd=8.28e+06u as=5.88e+11p ps=4.76e+06u
M1003 a_96_74# C VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR D a_96_74# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_96_74# A VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_257_74# B a_179_74# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.536e+11p ps=1.76e+06u
M1007 a_335_74# C a_257_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_96_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1009 a_179_74# A a_96_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
.ends

