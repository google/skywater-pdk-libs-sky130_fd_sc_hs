* File: sky130_fd_sc_hs__o32a_4.pxi.spice
* Created: Tue Sep  1 20:18:45 2020
* 
x_PM_SKY130_FD_SC_HS__O32A_4%A_83_256# N_A_83_256#_M1008_d N_A_83_256#_M1021_s
+ N_A_83_256#_M1004_d N_A_83_256#_M1003_d N_A_83_256#_c_161_n
+ N_A_83_256#_c_177_n N_A_83_256#_M1014_g N_A_83_256#_M1013_g
+ N_A_83_256#_c_163_n N_A_83_256#_c_164_n N_A_83_256#_c_179_n
+ N_A_83_256#_M1015_g N_A_83_256#_M1019_g N_A_83_256#_c_180_n
+ N_A_83_256#_M1016_g N_A_83_256#_M1024_g N_A_83_256#_c_181_n
+ N_A_83_256#_M1022_g N_A_83_256#_M1027_g N_A_83_256#_c_168_n
+ N_A_83_256#_c_169_n N_A_83_256#_c_170_n N_A_83_256#_c_171_n
+ N_A_83_256#_c_172_n N_A_83_256#_c_173_n N_A_83_256#_c_201_p
+ N_A_83_256#_c_174_n N_A_83_256#_c_184_n N_A_83_256#_c_233_p
+ N_A_83_256#_c_175_n PM_SKY130_FD_SC_HS__O32A_4%A_83_256#
x_PM_SKY130_FD_SC_HS__O32A_4%B1 N_B1_c_334_n N_B1_M1009_g N_B1_c_335_n
+ N_B1_c_336_n N_B1_c_337_n N_B1_c_338_n N_B1_M1008_g N_B1_c_339_n N_B1_c_340_n
+ N_B1_M1025_g N_B1_c_346_n N_B1_M1026_g N_B1_c_347_n N_B1_c_348_n N_B1_c_349_n
+ N_B1_c_341_n N_B1_c_350_n N_B1_c_351_n N_B1_c_453_p N_B1_c_352_n N_B1_c_353_n
+ N_B1_c_342_n N_B1_c_343_n B1 N_B1_c_344_n PM_SKY130_FD_SC_HS__O32A_4%B1
x_PM_SKY130_FD_SC_HS__O32A_4%B2 N_B2_c_490_n N_B2_M1004_g N_B2_c_491_n
+ N_B2_c_492_n N_B2_c_482_n N_B2_M1006_g N_B2_c_483_n N_B2_c_484_n N_B2_M1021_g
+ N_B2_c_485_n N_B2_c_486_n N_B2_M1023_g N_B2_c_487_n B2 N_B2_c_488_n
+ N_B2_c_489_n PM_SKY130_FD_SC_HS__O32A_4%B2
x_PM_SKY130_FD_SC_HS__O32A_4%A3 N_A3_M1000_g N_A3_c_562_n N_A3_c_568_n
+ N_A3_M1003_g N_A3_M1007_g N_A3_M1011_g N_A3_c_564_n N_A3_c_570_n A3
+ N_A3_c_566_n PM_SKY130_FD_SC_HS__O32A_4%A3
x_PM_SKY130_FD_SC_HS__O32A_4%A2 N_A2_c_634_n N_A2_M1010_g N_A2_c_626_n
+ N_A2_M1001_g N_A2_c_627_n N_A2_M1005_g N_A2_c_628_n N_A2_M1020_g N_A2_c_629_n
+ N_A2_c_630_n A2 A2 A2 A2 N_A2_c_632_n N_A2_c_652_n A2 N_A2_c_633_n
+ PM_SKY130_FD_SC_HS__O32A_4%A2
x_PM_SKY130_FD_SC_HS__O32A_4%A1 N_A1_c_725_n N_A1_M1017_g N_A1_c_726_n
+ N_A1_c_727_n N_A1_c_719_n N_A1_M1002_g N_A1_c_728_n N_A1_M1018_g N_A1_c_720_n
+ N_A1_c_721_n N_A1_M1012_g N_A1_c_722_n N_A1_c_729_n A1 N_A1_c_723_n
+ N_A1_c_724_n PM_SKY130_FD_SC_HS__O32A_4%A1
x_PM_SKY130_FD_SC_HS__O32A_4%VPWR N_VPWR_M1014_d N_VPWR_M1015_d N_VPWR_M1022_d
+ N_VPWR_M1026_d N_VPWR_M1017_d N_VPWR_c_789_n N_VPWR_c_790_n N_VPWR_c_791_n
+ N_VPWR_c_792_n N_VPWR_c_793_n N_VPWR_c_794_n N_VPWR_c_795_n N_VPWR_c_796_n
+ N_VPWR_c_797_n VPWR N_VPWR_c_798_n N_VPWR_c_799_n N_VPWR_c_800_n
+ N_VPWR_c_788_n N_VPWR_c_802_n N_VPWR_c_803_n N_VPWR_c_804_n
+ PM_SKY130_FD_SC_HS__O32A_4%VPWR
x_PM_SKY130_FD_SC_HS__O32A_4%X N_X_M1013_d N_X_M1024_d N_X_M1014_s N_X_M1016_s
+ N_X_c_886_n N_X_c_887_n N_X_c_888_n N_X_c_895_n N_X_c_889_n N_X_c_896_n
+ N_X_c_890_n N_X_c_897_n N_X_c_891_n N_X_c_892_n N_X_c_930_n X N_X_c_894_n
+ PM_SKY130_FD_SC_HS__O32A_4%X
x_PM_SKY130_FD_SC_HS__O32A_4%A_534_388# N_A_534_388#_M1009_s
+ N_A_534_388#_M1006_s N_A_534_388#_c_962_n
+ PM_SKY130_FD_SC_HS__O32A_4%A_534_388#
x_PM_SKY130_FD_SC_HS__O32A_4%A_961_392# N_A_961_392#_M1003_s
+ N_A_961_392#_M1007_s N_A_961_392#_M1020_s N_A_961_392#_c_980_n
+ N_A_961_392#_c_994_n N_A_961_392#_c_998_n N_A_961_392#_c_991_n
+ N_A_961_392#_c_981_n N_A_961_392#_c_982_n N_A_961_392#_c_983_n
+ PM_SKY130_FD_SC_HS__O32A_4%A_961_392#
x_PM_SKY130_FD_SC_HS__O32A_4%A_1234_392# N_A_1234_392#_M1010_d
+ N_A_1234_392#_M1018_s N_A_1234_392#_c_1031_n N_A_1234_392#_c_1038_n
+ N_A_1234_392#_c_1030_n N_A_1234_392#_c_1041_n
+ PM_SKY130_FD_SC_HS__O32A_4%A_1234_392#
x_PM_SKY130_FD_SC_HS__O32A_4%VGND N_VGND_M1013_s N_VGND_M1019_s N_VGND_M1027_s
+ N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1002_d N_VGND_c_1053_n N_VGND_c_1054_n
+ N_VGND_c_1055_n N_VGND_c_1056_n N_VGND_c_1057_n N_VGND_c_1058_n
+ N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n N_VGND_c_1062_n
+ N_VGND_c_1063_n N_VGND_c_1064_n N_VGND_c_1065_n N_VGND_c_1066_n VGND
+ N_VGND_c_1067_n N_VGND_c_1068_n N_VGND_c_1069_n N_VGND_c_1070_n
+ N_VGND_c_1071_n PM_SKY130_FD_SC_HS__O32A_4%VGND
x_PM_SKY130_FD_SC_HS__O32A_4%A_564_74# N_A_564_74#_M1008_s N_A_564_74#_M1025_s
+ N_A_564_74#_M1023_d N_A_564_74#_M1011_d N_A_564_74#_M1005_d
+ N_A_564_74#_M1012_s N_A_564_74#_c_1160_n N_A_564_74#_c_1161_n
+ N_A_564_74#_c_1162_n N_A_564_74#_c_1176_n N_A_564_74#_c_1163_n
+ N_A_564_74#_c_1164_n N_A_564_74#_c_1198_n N_A_564_74#_c_1165_n
+ N_A_564_74#_c_1208_n N_A_564_74#_c_1166_n N_A_564_74#_c_1167_n
+ N_A_564_74#_c_1168_n N_A_564_74#_c_1169_n N_A_564_74#_c_1204_n
+ N_A_564_74#_c_1217_n PM_SKY130_FD_SC_HS__O32A_4%A_564_74#
cc_1 VNB N_A_83_256#_c_161_n 0.0139124f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.675
cc_2 VNB N_A_83_256#_M1013_g 0.0224732f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.74
cc_3 VNB N_A_83_256#_c_163_n 0.00585843f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.355
cc_4 VNB N_A_83_256#_c_164_n 0.0110137f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.675
cc_5 VNB N_A_83_256#_M1019_g 0.0208918f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_6 VNB N_A_83_256#_M1024_g 0.0229607f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=0.74
cc_7 VNB N_A_83_256#_M1027_g 0.0231429f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=0.74
cc_8 VNB N_A_83_256#_c_168_n 0.013286f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.355
cc_9 VNB N_A_83_256#_c_169_n 0.00163584f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.445
cc_10 VNB N_A_83_256#_c_170_n 0.0915326f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.445
cc_11 VNB N_A_83_256#_c_171_n 0.0226784f $X=-0.19 $Y=-0.245 $X2=3.23 $Y2=1.195
cc_12 VNB N_A_83_256#_c_172_n 0.0013403f $X=-0.19 $Y=-0.245 $X2=3.395 $Y2=1.28
cc_13 VNB N_A_83_256#_c_173_n 0.00846832f $X=-0.19 $Y=-0.245 $X2=3.395 $Y2=1.92
cc_14 VNB N_A_83_256#_c_174_n 0.00267952f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=1.015
cc_15 VNB N_A_83_256#_c_175_n 0.00527666f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.195
cc_16 VNB N_B1_c_334_n 0.0219896f $X=-0.19 $Y=-0.245 $X2=3.255 $Y2=0.37
cc_17 VNB N_B1_c_335_n 0.013557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_336_n 0.016436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_337_n 0.0119858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_338_n 0.0189724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_339_n 0.020595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_340_n 0.0145703f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.43
cc_23 VNB N_B1_c_341_n 0.00530224f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.355
cc_24 VNB N_B1_c_342_n 0.00489941f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.765
cc_25 VNB N_B1_c_343_n 0.0213149f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_26 VNB N_B1_c_344_n 0.00267016f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_27 VNB N_B2_c_482_n 0.0141814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B2_c_483_n 0.0280227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B2_c_484_n 0.0151192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B2_c_485_n 0.0302534f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.675
cc_31 VNB N_B2_c_486_n 0.0158157f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_32 VNB N_B2_c_487_n 0.0110645f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.355
cc_33 VNB N_B2_c_488_n 0.0236629f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_34 VNB N_B2_c_489_n 9.04634e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_35 VNB N_A3_M1000_g 0.022736f $X=-0.19 $Y=-0.245 $X2=3.26 $Y2=1.94
cc_36 VNB N_A3_c_562_n 0.0084209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A3_M1011_g 0.0217763f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_38 VNB N_A3_c_564_n 0.00799726f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.74
cc_39 VNB A3 0.0124579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A3_c_566_n 0.044114f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.28
cc_41 VNB N_A2_c_626_n 0.0162939f $X=-0.19 $Y=-0.245 $X2=5.25 $Y2=1.96
cc_42 VNB N_A2_c_627_n 0.0156098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A2_c_628_n 0.023489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A2_c_629_n 0.029645f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_45 VNB N_A2_c_630_n 0.00499367f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_46 VNB A2 0.0116853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A2_c_632_n 0.0326934f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.28
cc_48 VNB N_A2_c_633_n 0.00960991f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_49 VNB N_A1_c_719_n 0.0172606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A1_c_720_n 0.0298031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A1_c_721_n 0.0223976f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.675
cc_52 VNB N_A1_c_722_n 0.00981662f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.28
cc_53 VNB N_A1_c_723_n 0.0352436f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.43
cc_54 VNB N_A1_c_724_n 0.0111425f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.675
cc_55 VNB N_VPWR_c_788_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_X_c_886_n 0.00341655f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.43
cc_57 VNB N_X_c_887_n 0.00221303f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_58 VNB N_X_c_888_n 0.00932569f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_59 VNB N_X_c_889_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.675
cc_60 VNB N_X_c_890_n 0.00162994f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.28
cc_61 VNB N_X_c_891_n 0.00282884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_X_c_892_n 0.00154309f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.4
cc_63 VNB X 0.00825292f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.445
cc_64 VNB N_X_c_894_n 0.011349f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_65 VNB N_VGND_c_1053_n 0.0144497f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.74
cc_66 VNB N_VGND_c_1054_n 0.0355428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1055_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.355
cc_68 VNB N_VGND_c_1056_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_69 VNB N_VGND_c_1057_n 0.011586f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_70 VNB N_VGND_c_1058_n 0.00867401f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_71 VNB N_VGND_c_1059_n 0.00508214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1060_n 0.00947287f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=1.28
cc_73 VNB N_VGND_c_1061_n 0.020287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1062_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.355
cc_75 VNB N_VGND_c_1063_n 0.0627424f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_76 VNB N_VGND_c_1064_n 0.00632279f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_77 VNB N_VGND_c_1065_n 0.0186748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1066_n 0.00613276f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.445
cc_79 VNB N_VGND_c_1067_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1068_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1069_n 0.436015f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.445
cc_82 VNB N_VGND_c_1070_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.43
cc_83 VNB N_VGND_c_1071_n 0.00737978f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.522
cc_84 VNB N_A_564_74#_c_1160_n 0.00465679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_564_74#_c_1161_n 0.00230691f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.355
cc_86 VNB N_A_564_74#_c_1162_n 0.00418558f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.43
cc_87 VNB N_A_564_74#_c_1163_n 0.00670648f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.28
cc_88 VNB N_A_564_74#_c_1164_n 0.00400232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_564_74#_c_1165_n 0.00256835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_564_74#_c_1166_n 0.00206225f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=0.74
cc_91 VNB N_A_564_74#_c_1167_n 0.0139705f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.355
cc_92 VNB N_A_564_74#_c_1168_n 0.0189752f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_93 VNB N_A_564_74#_c_1169_n 0.00220179f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.445
cc_94 VPB N_A_83_256#_c_161_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.675
cc_95 VPB N_A_83_256#_c_177_n 0.0258526f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_96 VPB N_A_83_256#_c_164_n 7.14638e-19 $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.675
cc_97 VPB N_A_83_256#_c_179_n 0.0207875f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_98 VPB N_A_83_256#_c_180_n 0.0158167f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_99 VPB N_A_83_256#_c_181_n 0.0170592f $X=-0.19 $Y=1.66 $X2=2.025 $Y2=1.765
cc_100 VPB N_A_83_256#_c_170_n 0.0149062f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.445
cc_101 VPB N_A_83_256#_c_173_n 0.0014396f $X=-0.19 $Y=1.66 $X2=3.395 $Y2=1.92
cc_102 VPB N_A_83_256#_c_184_n 0.00230942f $X=-0.19 $Y=1.66 $X2=5.4 $Y2=2.105
cc_103 VPB N_B1_c_334_n 0.038166f $X=-0.19 $Y=1.66 $X2=3.255 $Y2=0.37
cc_104 VPB N_B1_c_346_n 0.0142313f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_105 VPB N_B1_c_347_n 0.0376771f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_106 VPB N_B1_c_348_n 0.0132199f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_107 VPB N_B1_c_349_n 0.07095f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.355
cc_108 VPB N_B1_c_350_n 0.0027505f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.675
cc_109 VPB N_B1_c_351_n 0.00329833f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_110 VPB N_B1_c_352_n 0.0202558f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_111 VPB N_B1_c_353_n 0.00198471f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_112 VPB N_B1_c_342_n 0.00339195f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_113 VPB N_B1_c_343_n 0.013955f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_114 VPB N_B1_c_344_n 0.00123343f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.445
cc_115 VPB N_B2_c_490_n 0.0153275f $X=-0.19 $Y=1.66 $X2=3.255 $Y2=0.37
cc_116 VPB N_B2_c_491_n 0.0140178f $X=-0.19 $Y=1.66 $X2=5.25 $Y2=1.96
cc_117 VPB N_B2_c_492_n 0.0104353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_B2_c_482_n 0.0261945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_B2_c_489_n 0.00468087f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_120 VPB N_A3_c_562_n 0.00646578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A3_c_568_n 0.0220939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A3_c_564_n 0.00408276f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_123 VPB N_A3_c_570_n 0.0232861f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_124 VPB N_A2_c_634_n 0.0173854f $X=-0.19 $Y=1.66 $X2=3.255 $Y2=0.37
cc_125 VPB N_A2_c_628_n 0.0439634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A2_c_630_n 0.0238249f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_127 VPB A2 0.00227558f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.28
cc_128 VPB A2 0.00614495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A2_c_633_n 0.00476546f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.445
cc_130 VPB N_A1_c_725_n 0.0168203f $X=-0.19 $Y=1.66 $X2=3.255 $Y2=0.37
cc_131 VPB N_A1_c_726_n 0.00818126f $X=-0.19 $Y=1.66 $X2=5.25 $Y2=1.96
cc_132 VPB N_A1_c_727_n 0.0104445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A1_c_728_n 0.0154793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A1_c_729_n 0.0101608f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_135 VPB N_A1_c_723_n 0.00513583f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.43
cc_136 VPB N_VPWR_c_789_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_137 VPB N_VPWR_c_790_n 0.0570389f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.28
cc_138 VPB N_VPWR_c_791_n 0.00651803f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.43
cc_139 VPB N_VPWR_c_792_n 0.0190152f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_140 VPB N_VPWR_c_793_n 0.00724875f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_141 VPB N_VPWR_c_794_n 0.00517639f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.28
cc_142 VPB N_VPWR_c_795_n 0.00396467f $X=-0.19 $Y=1.66 $X2=2.025 $Y2=1.765
cc_143 VPB N_VPWR_c_796_n 0.0456519f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=1.28
cc_144 VPB N_VPWR_c_797_n 0.00510271f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=0.74
cc_145 VPB N_VPWR_c_798_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.562 $Y2=1.355
cc_146 VPB N_VPWR_c_799_n 0.0602951f $X=-0.19 $Y=1.66 $X2=3.395 $Y2=1.92
cc_147 VPB N_VPWR_c_800_n 0.0320405f $X=-0.19 $Y=1.66 $X2=5.4 $Y2=2.105
cc_148 VPB N_VPWR_c_788_n 0.0960468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_802_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_803_n 0.00614127f $X=-0.19 $Y=1.66 $X2=3.395 $Y2=1.015
cc_151 VPB N_VPWR_c_804_n 0.00601668f $X=-0.19 $Y=1.66 $X2=3.41 $Y2=2.095
cc_152 VPB N_X_c_895_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_153 VPB N_X_c_896_n 0.00618174f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_154 VPB N_X_c_897_n 0.00327585f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_155 VPB N_A_534_388#_c_962_n 0.00907611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_961_392#_c_980_n 0.0111223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_961_392#_c_981_n 0.0186878f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.355
cc_158 VPB N_A_961_392#_c_982_n 0.0188655f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_159 VPB N_A_961_392#_c_983_n 0.00704942f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_160 VPB N_A_1234_392#_c_1030_n 0.0026721f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=1.765
cc_161 N_A_83_256#_c_181_n N_B1_c_334_n 0.0168243f $X=2.025 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_83_256#_c_170_n N_B1_c_334_n 0.0138348f $X=2.1 $Y=1.445 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_83_256#_c_171_n N_B1_c_334_n 0.00541058f $X=3.23 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_83_256#_c_173_n N_B1_c_334_n 0.00128966f $X=3.395 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_83_256#_c_175_n N_B1_c_334_n 9.65797e-19 $X=2.27 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A_83_256#_c_170_n N_B1_c_335_n 0.00426339f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_167 N_A_83_256#_c_171_n N_B1_c_335_n 0.00402633f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_168 N_A_83_256#_c_173_n N_B1_c_335_n 0.005066f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_169 N_A_83_256#_c_175_n N_B1_c_335_n 0.00305315f $X=2.27 $Y=1.195 $X2=0 $Y2=0
cc_170 N_A_83_256#_c_171_n N_B1_c_336_n 0.00795139f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_171 N_A_83_256#_M1027_g N_B1_c_337_n 0.00426339f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_83_256#_c_171_n N_B1_c_337_n 0.00748939f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_173 N_A_83_256#_c_172_n N_B1_c_338_n 0.00255236f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_174 N_A_83_256#_c_172_n N_B1_c_339_n 0.0172734f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_175 N_A_83_256#_c_174_n N_B1_c_339_n 0.00201739f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_176 N_A_83_256#_c_172_n N_B1_c_340_n 0.00114575f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_177 N_A_83_256#_c_201_p N_B1_c_340_n 0.00559119f $X=3.395 $Y=0.81 $X2=0 $Y2=0
cc_178 N_A_83_256#_c_174_n N_B1_c_340_n 0.00713217f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_179 N_A_83_256#_c_173_n N_B1_c_346_n 7.2406e-19 $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_180 N_A_83_256#_c_184_n N_B1_c_346_n 0.010934f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_181 N_A_83_256#_c_184_n N_B1_c_349_n 0.0116343f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_182 N_A_83_256#_c_171_n N_B1_c_341_n 0.00724703f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_183 N_A_83_256#_c_172_n N_B1_c_341_n 0.0020413f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_184 N_A_83_256#_c_173_n N_B1_c_350_n 0.0170913f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_185 N_A_83_256#_M1004_d N_B1_c_351_n 0.00378224f $X=3.26 $Y=1.94 $X2=0 $Y2=0
cc_186 N_A_83_256#_M1003_d N_B1_c_351_n 0.00435327f $X=5.25 $Y=1.96 $X2=0 $Y2=0
cc_187 N_A_83_256#_c_173_n N_B1_c_351_n 0.0183569f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_188 N_A_83_256#_c_184_n N_B1_c_351_n 0.117556f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_189 N_A_83_256#_c_184_n N_B1_c_352_n 0.0476324f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_190 N_A_83_256#_c_174_n N_B1_c_342_n 0.00281519f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_191 N_A_83_256#_c_184_n N_B1_c_342_n 0.0252946f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_192 N_A_83_256#_c_184_n N_B1_c_343_n 0.00104009f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_193 N_A_83_256#_c_170_n N_B1_c_344_n 0.00104697f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_194 N_A_83_256#_c_171_n N_B1_c_344_n 0.0242401f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_195 N_A_83_256#_c_173_n N_B1_c_344_n 0.0141794f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_196 N_A_83_256#_c_175_n N_B1_c_344_n 0.0120085f $X=2.27 $Y=1.195 $X2=0 $Y2=0
cc_197 N_A_83_256#_c_173_n N_B2_c_490_n 0.0062287f $X=3.395 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_83_256#_c_173_n N_B2_c_491_n 0.0149534f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_199 N_A_83_256#_c_171_n N_B2_c_492_n 0.0023689f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_200 N_A_83_256#_c_173_n N_B2_c_492_n 0.00283456f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_201 N_A_83_256#_c_173_n N_B2_c_482_n 0.00936264f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_202 N_A_83_256#_c_174_n N_B2_c_482_n 0.00766854f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_203 N_A_83_256#_c_184_n N_B2_c_482_n 0.0116934f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_204 N_A_83_256#_c_184_n N_B2_c_483_n 0.00539085f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_205 N_A_83_256#_c_201_p N_B2_c_484_n 4.63525e-19 $X=3.395 $Y=0.81 $X2=0 $Y2=0
cc_206 N_A_83_256#_c_174_n N_B2_c_484_n 0.0101141f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_207 N_A_83_256#_c_174_n N_B2_c_485_n 0.0154786f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_208 N_A_83_256#_c_174_n N_B2_c_486_n 0.00371982f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_209 N_A_83_256#_c_233_p N_B2_c_486_n 0.00399613f $X=4.395 $Y=0.81 $X2=0 $Y2=0
cc_210 N_A_83_256#_c_172_n N_B2_c_487_n 8.09549e-19 $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_211 N_A_83_256#_c_174_n N_B2_c_487_n 0.00676917f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_212 N_A_83_256#_c_172_n N_B2_c_488_n 0.00127419f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_213 N_A_83_256#_c_173_n N_B2_c_488_n 0.00337625f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_214 N_A_83_256#_c_172_n N_B2_c_489_n 4.77843e-19 $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_215 N_A_83_256#_c_173_n N_B2_c_489_n 0.0228292f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_216 N_A_83_256#_c_174_n N_B2_c_489_n 0.0245197f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_217 N_A_83_256#_c_184_n N_B2_c_489_n 0.0171779f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_218 N_A_83_256#_c_174_n N_A3_M1000_g 4.24543e-19 $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_219 N_A_83_256#_c_184_n N_A3_c_568_n 0.00887154f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_220 N_A_83_256#_c_184_n N_VPWR_M1026_d 0.0133294f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_221 N_A_83_256#_c_177_n N_VPWR_c_790_n 0.0100916f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A_83_256#_c_179_n N_VPWR_c_791_n 0.00777421f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_A_83_256#_c_180_n N_VPWR_c_791_n 0.0142149f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_224 N_A_83_256#_c_181_n N_VPWR_c_791_n 6.69644e-19 $X=2.025 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_A_83_256#_c_180_n N_VPWR_c_792_n 0.00413917f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_A_83_256#_c_181_n N_VPWR_c_792_n 0.00413917f $X=2.025 $Y=1.765 $X2=0
+ $Y2=0
cc_227 N_A_83_256#_c_180_n N_VPWR_c_793_n 7.24688e-19 $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A_83_256#_c_181_n N_VPWR_c_793_n 0.0150251f $X=2.025 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A_83_256#_c_169_n N_VPWR_c_793_n 0.00320315f $X=2.185 $Y=1.445 $X2=0
+ $Y2=0
cc_230 N_A_83_256#_c_170_n N_VPWR_c_793_n 0.00213758f $X=2.1 $Y=1.445 $X2=0
+ $Y2=0
cc_231 N_A_83_256#_c_171_n N_VPWR_c_793_n 0.00179271f $X=3.23 $Y=1.195 $X2=0
+ $Y2=0
cc_232 N_A_83_256#_c_175_n N_VPWR_c_793_n 0.00880609f $X=2.27 $Y=1.195 $X2=0
+ $Y2=0
cc_233 N_A_83_256#_c_177_n N_VPWR_c_798_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A_83_256#_c_179_n N_VPWR_c_798_n 0.00445602f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_A_83_256#_c_177_n N_VPWR_c_788_n 0.00861084f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A_83_256#_c_179_n N_VPWR_c_788_n 0.00857378f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A_83_256#_c_180_n N_VPWR_c_788_n 0.00818763f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_83_256#_c_181_n N_VPWR_c_788_n 0.00818763f $X=2.025 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A_83_256#_M1013_g N_X_c_886_n 0.0109683f $X=0.635 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_83_256#_c_168_n N_X_c_886_n 0.00709161f $X=0.562 $Y=1.355 $X2=0 $Y2=0
cc_241 N_A_83_256#_c_161_n N_X_c_887_n 0.0149993f $X=0.505 $Y=1.675 $X2=0 $Y2=0
cc_242 N_A_83_256#_c_177_n N_X_c_895_n 0.0120721f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_83_256#_c_179_n N_X_c_895_n 0.0124759f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_244 N_A_83_256#_c_180_n N_X_c_895_n 2.70252e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_83_256#_M1013_g N_X_c_889_n 0.00746201f $X=0.635 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A_83_256#_M1019_g N_X_c_889_n 0.00896067f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_83_256#_M1024_g N_X_c_889_n 6.1951e-19 $X=1.635 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A_83_256#_c_179_n N_X_c_896_n 0.0152224f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_83_256#_c_180_n N_X_c_896_n 0.0154193f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A_83_256#_c_181_n N_X_c_896_n 0.00263207f $X=2.025 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A_83_256#_c_169_n N_X_c_896_n 0.050529f $X=2.185 $Y=1.445 $X2=0 $Y2=0
cc_252 N_A_83_256#_c_170_n N_X_c_896_n 0.0176477f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_253 N_A_83_256#_M1019_g N_X_c_890_n 0.0143019f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_83_256#_M1024_g N_X_c_890_n 0.0126012f $X=1.635 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_83_256#_M1027_g N_X_c_890_n 0.00533726f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_83_256#_c_169_n N_X_c_890_n 0.0539257f $X=2.185 $Y=1.445 $X2=0 $Y2=0
cc_257 N_A_83_256#_c_170_n N_X_c_890_n 0.0110961f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_258 N_A_83_256#_c_180_n N_X_c_897_n 0.00644771f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A_83_256#_c_181_n N_X_c_897_n 0.00619894f $X=2.025 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A_83_256#_M1019_g N_X_c_891_n 6.14947e-19 $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_83_256#_M1024_g N_X_c_891_n 0.00878544f $X=1.635 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_83_256#_M1027_g N_X_c_891_n 0.00535397f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_83_256#_c_161_n N_X_c_892_n 0.00467185f $X=0.505 $Y=1.675 $X2=0 $Y2=0
cc_264 N_A_83_256#_c_177_n N_X_c_892_n 0.0100229f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A_83_256#_c_164_n N_X_c_892_n 0.00581793f $X=0.955 $Y=1.675 $X2=0 $Y2=0
cc_266 N_A_83_256#_c_179_n N_X_c_892_n 0.00513713f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A_83_256#_c_180_n N_X_c_892_n 6.04667e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A_83_256#_c_168_n N_X_c_892_n 0.0028273f $X=0.562 $Y=1.355 $X2=0 $Y2=0
cc_269 N_A_83_256#_c_169_n N_X_c_892_n 0.00562369f $X=2.185 $Y=1.445 $X2=0 $Y2=0
cc_270 N_A_83_256#_c_170_n N_X_c_892_n 8.53025e-19 $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_271 N_A_83_256#_M1013_g N_X_c_930_n 0.0104872f $X=0.635 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A_83_256#_c_163_n N_X_c_930_n 0.00361547f $X=0.865 $Y=1.355 $X2=0 $Y2=0
cc_273 N_A_83_256#_M1019_g N_X_c_930_n 0.00636589f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_83_256#_M1024_g N_X_c_930_n 8.53592e-19 $X=1.635 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A_83_256#_c_168_n N_X_c_930_n 3.57967e-19 $X=0.562 $Y=1.355 $X2=0 $Y2=0
cc_276 N_A_83_256#_c_169_n N_X_c_930_n 0.00175494f $X=2.185 $Y=1.445 $X2=0 $Y2=0
cc_277 N_A_83_256#_c_170_n N_X_c_930_n 0.00486665f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_278 N_A_83_256#_c_168_n X 0.00776373f $X=0.562 $Y=1.355 $X2=0 $Y2=0
cc_279 N_A_83_256#_c_184_n N_A_534_388#_M1006_s 0.00454772f $X=5.4 $Y=2.105
+ $X2=0 $Y2=0
cc_280 N_A_83_256#_M1004_d N_A_534_388#_c_962_n 0.00200816f $X=3.26 $Y=1.94
+ $X2=0 $Y2=0
cc_281 N_A_83_256#_c_184_n N_A_961_392#_M1003_s 0.00511055f $X=5.4 $Y=2.105
+ $X2=-0.19 $Y2=-0.245
cc_282 N_A_83_256#_M1003_d N_A_961_392#_c_980_n 0.00222916f $X=5.25 $Y=1.96
+ $X2=0 $Y2=0
cc_283 N_A_83_256#_c_175_n N_VGND_M1027_s 9.75702e-19 $X=2.27 $Y=1.195 $X2=0
+ $Y2=0
cc_284 N_A_83_256#_M1013_g N_VGND_c_1054_n 0.0153292f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_83_256#_c_168_n N_VGND_c_1054_n 5.27843e-19 $X=0.562 $Y=1.355 $X2=0
+ $Y2=0
cc_286 N_A_83_256#_M1013_g N_VGND_c_1055_n 0.00434272f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_83_256#_M1019_g N_VGND_c_1055_n 0.00434272f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_288 N_A_83_256#_M1019_g N_VGND_c_1056_n 0.00441895f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_83_256#_M1024_g N_VGND_c_1056_n 0.00580088f $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_290 N_A_83_256#_M1024_g N_VGND_c_1057_n 7.01214e-19 $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_291 N_A_83_256#_M1027_g N_VGND_c_1057_n 0.0125112f $X=2.19 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_83_256#_c_171_n N_VGND_c_1057_n 0.0177292f $X=3.23 $Y=1.195 $X2=0
+ $Y2=0
cc_293 N_A_83_256#_c_175_n N_VGND_c_1057_n 0.00721878f $X=2.27 $Y=1.195 $X2=0
+ $Y2=0
cc_294 N_A_83_256#_M1024_g N_VGND_c_1061_n 0.00434272f $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_295 N_A_83_256#_M1027_g N_VGND_c_1061_n 0.00383152f $X=2.19 $Y=0.74 $X2=0
+ $Y2=0
cc_296 N_A_83_256#_M1013_g N_VGND_c_1069_n 0.00824109f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_297 N_A_83_256#_M1019_g N_VGND_c_1069_n 0.00821294f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_298 N_A_83_256#_M1024_g N_VGND_c_1069_n 0.0082241f $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_83_256#_M1027_g N_VGND_c_1069_n 0.00758657f $X=2.19 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_83_256#_c_174_n N_A_564_74#_M1025_s 0.00250873f $X=4.23 $Y=1.015
+ $X2=0 $Y2=0
cc_301 N_A_83_256#_c_171_n N_A_564_74#_c_1160_n 0.0232013f $X=3.23 $Y=1.195
+ $X2=0 $Y2=0
cc_302 N_A_83_256#_M1008_d N_A_564_74#_c_1161_n 0.00168861f $X=3.255 $Y=0.37
+ $X2=0 $Y2=0
cc_303 N_A_83_256#_c_201_p N_A_564_74#_c_1161_n 0.0143448f $X=3.395 $Y=0.81
+ $X2=0 $Y2=0
cc_304 N_A_83_256#_c_174_n N_A_564_74#_c_1161_n 0.00347117f $X=4.23 $Y=1.015
+ $X2=0 $Y2=0
cc_305 N_A_83_256#_M1027_g N_A_564_74#_c_1162_n 6.04331e-19 $X=2.19 $Y=0.74
+ $X2=0 $Y2=0
cc_306 N_A_83_256#_c_174_n N_A_564_74#_c_1176_n 0.0204865f $X=4.23 $Y=1.015
+ $X2=0 $Y2=0
cc_307 N_A_83_256#_M1021_s N_A_564_74#_c_1163_n 0.00237953f $X=4.185 $Y=0.37
+ $X2=0 $Y2=0
cc_308 N_A_83_256#_c_174_n N_A_564_74#_c_1163_n 0.00347117f $X=4.23 $Y=1.015
+ $X2=0 $Y2=0
cc_309 N_A_83_256#_c_233_p N_A_564_74#_c_1163_n 0.0192294f $X=4.395 $Y=0.81
+ $X2=0 $Y2=0
cc_310 N_B1_c_334_n N_B2_c_490_n 0.0271284f $X=2.595 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_311 N_B1_c_350_n N_B2_c_490_n 0.00598861f $X=2.77 $Y=2.36 $X2=-0.19
+ $Y2=-0.245
cc_312 N_B1_c_351_n N_B2_c_490_n 0.0146379f $X=5.735 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_313 N_B1_c_341_n N_B2_c_491_n 0.00348858f $X=3.18 $Y=1.165 $X2=0 $Y2=0
cc_314 N_B1_c_351_n N_B2_c_491_n 4.2495e-19 $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_315 N_B1_c_334_n N_B2_c_492_n 0.00564384f $X=2.595 $Y=1.865 $X2=0 $Y2=0
cc_316 N_B1_c_336_n N_B2_c_492_n 0.00348858f $X=3.105 $Y=1.165 $X2=0 $Y2=0
cc_317 N_B1_c_350_n N_B2_c_492_n 8.12804e-19 $X=2.77 $Y=2.36 $X2=0 $Y2=0
cc_318 N_B1_c_344_n N_B2_c_492_n 2.86983e-19 $X=2.77 $Y=1.615 $X2=0 $Y2=0
cc_319 N_B1_c_334_n N_B2_c_482_n 0.00236341f $X=2.595 $Y=1.865 $X2=0 $Y2=0
cc_320 N_B1_c_339_n N_B2_c_482_n 0.0120559f $X=3.535 $Y=1.165 $X2=0 $Y2=0
cc_321 N_B1_c_346_n N_B2_c_482_n 0.0378279f $X=4.085 $Y=3.015 $X2=0 $Y2=0
cc_322 N_B1_c_348_n N_B2_c_482_n 0.00286983f $X=4.16 $Y=3.09 $X2=0 $Y2=0
cc_323 N_B1_c_351_n N_B2_c_482_n 0.0106731f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_324 N_B1_c_346_n N_B2_c_483_n 0.00983426f $X=4.085 $Y=3.015 $X2=0 $Y2=0
cc_325 N_B1_c_342_n N_B2_c_483_n 6.33942e-19 $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_326 N_B1_c_343_n N_B2_c_483_n 0.00821351f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_327 N_B1_c_340_n N_B2_c_484_n 0.0203621f $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_328 N_B1_c_342_n N_B2_c_485_n 0.00123953f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_329 N_B1_c_343_n N_B2_c_485_n 0.0126816f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_330 N_B1_c_339_n N_B2_c_487_n 0.0100546f $X=3.535 $Y=1.165 $X2=0 $Y2=0
cc_331 N_B1_c_346_n N_B2_c_489_n 0.00150864f $X=4.085 $Y=3.015 $X2=0 $Y2=0
cc_332 N_B1_c_342_n N_B2_c_489_n 0.0195613f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_333 N_B1_c_343_n N_B2_c_489_n 0.00447962f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_334 N_B1_c_349_n N_A3_c_562_n 0.00373034f $X=4.655 $Y=3.015 $X2=0 $Y2=0
cc_335 N_B1_c_352_n N_A3_c_562_n 0.00707722f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_336 N_B1_c_342_n N_A3_c_562_n 0.00122954f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_337 N_B1_c_343_n N_A3_c_562_n 0.0137874f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_338 N_B1_c_349_n N_A3_c_568_n 0.0352038f $X=4.655 $Y=3.015 $X2=0 $Y2=0
cc_339 N_B1_c_351_n N_A3_c_568_n 0.0110921f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_340 N_B1_c_352_n N_A3_c_568_n 0.00443784f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_341 N_B1_c_352_n N_A3_c_564_n 0.00442139f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_342 N_B1_c_351_n N_A3_c_570_n 0.0117565f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_343 N_B1_c_352_n N_A3_c_570_n 0.00762892f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_344 N_B1_c_353_n N_A3_c_570_n 0.0046977f $X=5.82 $Y=2.36 $X2=0 $Y2=0
cc_345 N_B1_c_352_n A3 0.0490884f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_346 N_B1_c_342_n A3 0.0035661f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_347 N_B1_c_343_n A3 2.16867e-19 $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_348 N_B1_c_352_n N_A3_c_566_n 0.00366609f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_349 N_B1_c_343_n N_A3_c_566_n 0.00323048f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_350 N_B1_c_351_n N_A2_c_634_n 0.00191892f $X=5.735 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_351 N_B1_c_353_n N_A2_c_634_n 0.00689562f $X=5.82 $Y=2.36 $X2=-0.19
+ $Y2=-0.245
cc_352 N_B1_c_352_n N_A2_c_630_n 0.00247751f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_353 N_B1_c_353_n N_A2_c_630_n 7.7174e-19 $X=5.82 $Y=2.36 $X2=0 $Y2=0
cc_354 N_B1_c_352_n A2 0.0106093f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_355 N_B1_c_351_n N_VPWR_M1026_d 0.00633878f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_356 N_B1_c_334_n N_VPWR_c_793_n 0.0157391f $X=2.595 $Y=1.865 $X2=0 $Y2=0
cc_357 N_B1_c_346_n N_VPWR_c_794_n 0.00331738f $X=4.085 $Y=3.015 $X2=0 $Y2=0
cc_358 N_B1_c_347_n N_VPWR_c_794_n 0.022065f $X=4.58 $Y=3.09 $X2=0 $Y2=0
cc_359 N_B1_c_349_n N_VPWR_c_794_n 0.00403053f $X=4.655 $Y=3.015 $X2=0 $Y2=0
cc_360 N_B1_c_351_n N_VPWR_c_794_n 0.0245011f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_361 N_B1_c_334_n N_VPWR_c_796_n 0.00547215f $X=2.595 $Y=1.865 $X2=0 $Y2=0
cc_362 N_B1_c_348_n N_VPWR_c_796_n 0.00656219f $X=4.16 $Y=3.09 $X2=0 $Y2=0
cc_363 N_B1_c_347_n N_VPWR_c_799_n 0.00716255f $X=4.58 $Y=3.09 $X2=0 $Y2=0
cc_364 N_B1_c_334_n N_VPWR_c_788_n 0.00539454f $X=2.595 $Y=1.865 $X2=0 $Y2=0
cc_365 N_B1_c_347_n N_VPWR_c_788_n 0.00856279f $X=4.58 $Y=3.09 $X2=0 $Y2=0
cc_366 N_B1_c_348_n N_VPWR_c_788_n 0.00622128f $X=4.16 $Y=3.09 $X2=0 $Y2=0
cc_367 N_B1_c_351_n N_VPWR_c_788_n 0.0171185f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_368 N_B1_c_350_n N_A_534_388#_M1009_s 0.00790577f $X=2.77 $Y=2.36 $X2=-0.19
+ $Y2=-0.245
cc_369 N_B1_c_351_n N_A_534_388#_M1009_s 0.0102686f $X=5.735 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_370 N_B1_c_453_p N_A_534_388#_M1009_s 0.0025282f $X=2.855 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_371 N_B1_c_351_n N_A_534_388#_M1006_s 0.00393062f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_372 N_B1_c_334_n N_A_534_388#_c_962_n 0.00800586f $X=2.595 $Y=1.865 $X2=0
+ $Y2=0
cc_373 N_B1_c_346_n N_A_534_388#_c_962_n 0.00310189f $X=4.085 $Y=3.015 $X2=0
+ $Y2=0
cc_374 N_B1_c_348_n N_A_534_388#_c_962_n 3.60338e-19 $X=4.16 $Y=3.09 $X2=0 $Y2=0
cc_375 N_B1_c_351_n N_A_534_388#_c_962_n 0.0629112f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_376 N_B1_c_453_p N_A_534_388#_c_962_n 0.0103504f $X=2.855 $Y=2.445 $X2=0
+ $Y2=0
cc_377 N_B1_c_351_n N_A_961_392#_M1003_s 0.00509354f $X=5.735 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_378 N_B1_c_351_n N_A_961_392#_M1007_s 0.00298057f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_379 N_B1_c_353_n N_A_961_392#_M1007_s 0.0051458f $X=5.82 $Y=2.36 $X2=0 $Y2=0
cc_380 N_B1_c_349_n N_A_961_392#_c_980_n 0.00306725f $X=4.655 $Y=3.015 $X2=0
+ $Y2=0
cc_381 N_B1_c_351_n N_A_961_392#_c_980_n 0.064978f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_382 N_B1_c_351_n N_A_961_392#_c_991_n 0.0122365f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_383 N_B1_c_353_n N_A_1234_392#_c_1031_n 0.0144376f $X=5.82 $Y=2.36 $X2=0
+ $Y2=0
cc_384 N_B1_c_338_n N_VGND_c_1057_n 0.00176715f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_385 N_B1_c_338_n N_VGND_c_1063_n 0.00278247f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_386 N_B1_c_340_n N_VGND_c_1063_n 0.00278271f $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_387 N_B1_c_338_n N_VGND_c_1069_n 0.00358425f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_388 N_B1_c_340_n N_VGND_c_1069_n 0.0035414f $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_389 N_B1_c_337_n N_A_564_74#_c_1160_n 0.00638349f $X=2.855 $Y=1.165 $X2=0
+ $Y2=0
cc_390 N_B1_c_338_n N_A_564_74#_c_1160_n 0.00694622f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_391 N_B1_c_340_n N_A_564_74#_c_1160_n 6.20636e-19 $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_392 N_B1_c_338_n N_A_564_74#_c_1161_n 0.0100711f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_393 N_B1_c_339_n N_A_564_74#_c_1161_n 2.67777e-19 $X=3.535 $Y=1.165 $X2=0
+ $Y2=0
cc_394 N_B1_c_340_n N_A_564_74#_c_1161_n 0.0109066f $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_395 N_B1_c_338_n N_A_564_74#_c_1162_n 0.00281658f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_396 N_B1_c_352_n N_A_564_74#_c_1164_n 0.0063124f $X=5.735 $Y=1.765 $X2=0
+ $Y2=0
cc_397 N_B1_c_342_n N_A_564_74#_c_1164_n 0.00351334f $X=4.66 $Y=1.615 $X2=0
+ $Y2=0
cc_398 N_B1_c_343_n N_A_564_74#_c_1164_n 5.96818e-19 $X=4.66 $Y=1.615 $X2=0
+ $Y2=0
cc_399 N_B2_c_486_n N_A3_M1000_g 0.00961692f $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_400 N_B2_c_485_n A3 4.16793e-19 $X=4.535 $Y=1.165 $X2=0 $Y2=0
cc_401 N_B2_c_485_n N_A3_c_566_n 0.00961692f $X=4.535 $Y=1.165 $X2=0 $Y2=0
cc_402 N_B2_c_482_n N_VPWR_c_794_n 2.33869e-19 $X=3.635 $Y=1.865 $X2=0 $Y2=0
cc_403 N_B2_c_490_n N_VPWR_c_796_n 0.00401361f $X=3.185 $Y=1.865 $X2=0 $Y2=0
cc_404 N_B2_c_482_n N_VPWR_c_796_n 0.00401361f $X=3.635 $Y=1.865 $X2=0 $Y2=0
cc_405 N_B2_c_490_n N_VPWR_c_788_n 0.00539454f $X=3.185 $Y=1.865 $X2=0 $Y2=0
cc_406 N_B2_c_482_n N_VPWR_c_788_n 0.00539454f $X=3.635 $Y=1.865 $X2=0 $Y2=0
cc_407 N_B2_c_490_n N_A_534_388#_c_962_n 0.0147454f $X=3.185 $Y=1.865 $X2=0
+ $Y2=0
cc_408 N_B2_c_482_n N_A_534_388#_c_962_n 0.010745f $X=3.635 $Y=1.865 $X2=0 $Y2=0
cc_409 N_B2_c_484_n N_VGND_c_1063_n 0.00278247f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_410 N_B2_c_486_n N_VGND_c_1063_n 0.00278271f $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_411 N_B2_c_484_n N_VGND_c_1069_n 0.00354796f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_412 N_B2_c_486_n N_VGND_c_1069_n 0.00355038f $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_413 N_B2_c_484_n N_A_564_74#_c_1176_n 0.00539089f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_414 N_B2_c_486_n N_A_564_74#_c_1176_n 5.81199e-19 $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_415 N_B2_c_487_n N_A_564_74#_c_1176_n 4.55305e-19 $X=4.09 $Y=1.165 $X2=0
+ $Y2=0
cc_416 N_B2_c_484_n N_A_564_74#_c_1163_n 0.00806723f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_417 N_B2_c_485_n N_A_564_74#_c_1163_n 4.55221e-19 $X=4.535 $Y=1.165 $X2=0
+ $Y2=0
cc_418 N_B2_c_486_n N_A_564_74#_c_1163_n 0.0137079f $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_419 N_B2_c_484_n N_A_564_74#_c_1169_n 0.00253515f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_420 N_A3_c_570_n N_A2_c_634_n 0.0305207f $X=5.652 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_421 N_A3_M1011_g N_A2_c_626_n 0.0110549f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_422 N_A3_M1011_g N_A2_c_629_n 0.0119082f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_423 A3 N_A2_c_629_n 0.00137288f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_424 N_A3_c_564_n N_A2_c_630_n 0.0119082f $X=5.652 $Y=1.75 $X2=0 $Y2=0
cc_425 N_A3_c_564_n A2 6.38729e-19 $X=5.652 $Y=1.75 $X2=0 $Y2=0
cc_426 N_A3_c_566_n N_A2_c_632_n 0.0119082f $X=5.66 $Y=1.345 $X2=0 $Y2=0
cc_427 N_A3_M1011_g N_A2_c_652_n 2.7656e-19 $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_428 A3 N_A2_c_652_n 0.0149466f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_429 N_A3_c_566_n N_A2_c_652_n 7.57327e-19 $X=5.66 $Y=1.345 $X2=0 $Y2=0
cc_430 N_A3_c_568_n N_VPWR_c_794_n 3.15949e-19 $X=5.175 $Y=1.885 $X2=0 $Y2=0
cc_431 N_A3_c_568_n N_VPWR_c_799_n 0.00291649f $X=5.175 $Y=1.885 $X2=0 $Y2=0
cc_432 N_A3_c_570_n N_VPWR_c_799_n 0.00291649f $X=5.652 $Y=1.885 $X2=0 $Y2=0
cc_433 N_A3_c_568_n N_VPWR_c_788_n 0.00360381f $X=5.175 $Y=1.885 $X2=0 $Y2=0
cc_434 N_A3_c_570_n N_VPWR_c_788_n 0.00359789f $X=5.652 $Y=1.885 $X2=0 $Y2=0
cc_435 N_A3_c_568_n N_A_961_392#_c_980_n 0.0114055f $X=5.175 $Y=1.885 $X2=0
+ $Y2=0
cc_436 N_A3_c_570_n N_A_961_392#_c_980_n 0.0114016f $X=5.652 $Y=1.885 $X2=0
+ $Y2=0
cc_437 N_A3_c_570_n N_A_961_392#_c_994_n 5.34839e-19 $X=5.652 $Y=1.885 $X2=0
+ $Y2=0
cc_438 N_A3_c_570_n N_A_961_392#_c_991_n 2.88318e-19 $X=5.652 $Y=1.885 $X2=0
+ $Y2=0
cc_439 N_A3_M1000_g N_VGND_c_1058_n 0.00148871f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_440 N_A3_M1011_g N_VGND_c_1058_n 0.00198878f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_441 N_A3_M1000_g N_VGND_c_1063_n 0.00461464f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_442 N_A3_M1011_g N_VGND_c_1065_n 0.00456932f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_443 N_A3_M1000_g N_VGND_c_1069_n 0.00451999f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_444 N_A3_M1011_g N_VGND_c_1069_n 0.00443718f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_445 N_A3_M1000_g N_A_564_74#_c_1163_n 0.00118927f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_446 N_A3_M1000_g N_A_564_74#_c_1198_n 0.0104635f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_447 N_A3_M1011_g N_A_564_74#_c_1198_n 0.0101963f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_448 A3 N_A_564_74#_c_1198_n 0.036068f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_449 N_A3_c_566_n N_A_564_74#_c_1198_n 0.00430721f $X=5.66 $Y=1.345 $X2=0
+ $Y2=0
cc_450 N_A3_M1000_g N_A_564_74#_c_1165_n 3.11133e-19 $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_451 N_A3_M1011_g N_A_564_74#_c_1165_n 0.00560871f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_452 N_A3_M1011_g N_A_564_74#_c_1204_n 2.51849e-19 $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_453 A3 N_A_564_74#_c_1204_n 2.88494e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_454 N_A2_c_634_n N_A1_c_725_n 0.0270293f $X=6.095 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_455 N_A2_c_633_n N_A1_c_726_n 0.00514608f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_456 N_A2_c_629_n N_A1_c_727_n 8.16592e-19 $X=6.205 $Y=1.235 $X2=0 $Y2=0
cc_457 N_A2_c_630_n N_A1_c_727_n 0.00674971f $X=6.205 $Y=1.6 $X2=0 $Y2=0
cc_458 N_A2_c_633_n N_A1_c_727_n 0.00610695f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_459 N_A2_c_627_n N_A1_c_719_n 0.00828772f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_460 N_A2_c_628_n N_A1_c_728_n 0.035278f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_461 N_A2_c_628_n N_A1_c_720_n 0.0125022f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_462 A2 N_A1_c_720_n 8.24499e-19 $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_463 N_A2_c_633_n N_A1_c_720_n 0.00558949f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_464 N_A2_c_629_n N_A1_c_722_n 0.00828772f $X=6.205 $Y=1.235 $X2=0 $Y2=0
cc_465 N_A2_c_632_n N_A1_c_722_n 0.00478184f $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_466 N_A2_c_652_n N_A1_c_722_n 2.55438e-19 $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_467 N_A2_c_633_n N_A1_c_729_n 0.00612479f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_468 N_A2_c_628_n N_A1_c_723_n 0.021792f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_469 N_A2_c_630_n N_A1_c_723_n 0.00478184f $X=6.205 $Y=1.6 $X2=0 $Y2=0
cc_470 A2 N_A1_c_723_n 8.80533e-19 $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_471 N_A2_c_652_n N_A1_c_723_n 9.78829e-19 $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_472 N_A2_c_633_n N_A1_c_723_n 0.0139494f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_473 N_A2_c_629_n N_A1_c_724_n 0.00142867f $X=6.205 $Y=1.235 $X2=0 $Y2=0
cc_474 N_A2_c_632_n N_A1_c_724_n 0.00149364f $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_475 N_A2_c_652_n N_A1_c_724_n 0.0111493f $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_476 N_A2_c_633_n N_A1_c_724_n 0.0331366f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_477 N_A2_c_634_n N_VPWR_c_795_n 7.02217e-19 $X=6.095 $Y=1.885 $X2=0 $Y2=0
cc_478 N_A2_c_628_n N_VPWR_c_795_n 0.00125269f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_479 N_A2_c_634_n N_VPWR_c_799_n 0.00291563f $X=6.095 $Y=1.885 $X2=0 $Y2=0
cc_480 N_A2_c_628_n N_VPWR_c_800_n 0.00445602f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_481 N_A2_c_634_n N_VPWR_c_788_n 0.00361064f $X=6.095 $Y=1.885 $X2=0 $Y2=0
cc_482 N_A2_c_628_n N_VPWR_c_788_n 0.00441311f $X=7.655 $Y=1.885 $X2=0 $Y2=0
cc_483 N_A2_c_634_n N_A_961_392#_c_980_n 0.0106844f $X=6.095 $Y=1.885 $X2=0
+ $Y2=0
cc_484 N_A2_c_634_n N_A_961_392#_c_994_n 0.00442991f $X=6.095 $Y=1.885 $X2=0
+ $Y2=0
cc_485 N_A2_c_628_n N_A_961_392#_c_998_n 0.0105677f $X=7.655 $Y=1.885 $X2=0
+ $Y2=0
cc_486 A2 N_A_961_392#_c_998_n 0.00296232f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_487 N_A2_c_634_n N_A_961_392#_c_991_n 0.00829944f $X=6.095 $Y=1.885 $X2=0
+ $Y2=0
cc_488 A2 N_A_961_392#_c_991_n 0.00237965f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_489 N_A2_c_628_n N_A_961_392#_c_981_n 0.00795639f $X=7.655 $Y=1.885 $X2=0
+ $Y2=0
cc_490 N_A2_c_628_n N_A_961_392#_c_982_n 0.00324938f $X=7.655 $Y=1.885 $X2=0
+ $Y2=0
cc_491 A2 N_A_961_392#_c_982_n 0.0232636f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_492 N_A2_c_628_n N_A_961_392#_c_983_n 6.02976e-19 $X=7.655 $Y=1.885 $X2=0
+ $Y2=0
cc_493 A2 N_A_961_392#_c_983_n 8.52067e-19 $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_494 N_A2_c_634_n N_A_1234_392#_c_1031_n 0.0075608f $X=6.095 $Y=1.885 $X2=0
+ $Y2=0
cc_495 N_A2_c_630_n N_A_1234_392#_c_1031_n 0.00147472f $X=6.205 $Y=1.6 $X2=0
+ $Y2=0
cc_496 A2 N_A_1234_392#_c_1031_n 0.017928f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_497 N_A2_c_633_n N_A_1234_392#_c_1031_n 0.0515565f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_498 N_A2_c_628_n N_A_1234_392#_c_1030_n 0.00340355f $X=7.655 $Y=1.885 $X2=0
+ $Y2=0
cc_499 N_A2_c_633_n N_A_1234_392#_c_1030_n 0.0256037f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_500 N_A2_c_626_n N_VGND_c_1059_n 0.00312943f $X=6.11 $Y=1.085 $X2=0 $Y2=0
cc_501 N_A2_c_627_n N_VGND_c_1059_n 0.0070913f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_502 N_A2_c_626_n N_VGND_c_1065_n 0.00434272f $X=6.11 $Y=1.085 $X2=0 $Y2=0
cc_503 N_A2_c_627_n N_VGND_c_1067_n 0.00383152f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_504 N_A2_c_626_n N_VGND_c_1069_n 0.00433282f $X=6.11 $Y=1.085 $X2=0 $Y2=0
cc_505 N_A2_c_627_n N_VGND_c_1069_n 0.0037147f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_506 N_A2_c_626_n N_A_564_74#_c_1165_n 0.00639171f $X=6.11 $Y=1.085 $X2=0
+ $Y2=0
cc_507 N_A2_c_627_n N_A_564_74#_c_1165_n 6.25537e-19 $X=6.61 $Y=1.085 $X2=0
+ $Y2=0
cc_508 N_A2_c_626_n N_A_564_74#_c_1208_n 0.00925007f $X=6.11 $Y=1.085 $X2=0
+ $Y2=0
cc_509 N_A2_c_627_n N_A_564_74#_c_1208_n 0.0111557f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_510 N_A2_c_629_n N_A_564_74#_c_1208_n 0.00458615f $X=6.205 $Y=1.235 $X2=0
+ $Y2=0
cc_511 N_A2_c_652_n N_A_564_74#_c_1208_n 0.0223703f $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_512 N_A2_c_633_n N_A_564_74#_c_1208_n 0.00783756f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_513 N_A2_c_628_n N_A_564_74#_c_1167_n 0.00347477f $X=7.655 $Y=1.885 $X2=0
+ $Y2=0
cc_514 A2 N_A_564_74#_c_1167_n 0.0183141f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_515 N_A2_c_633_n N_A_564_74#_c_1167_n 0.00735461f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_516 N_A2_c_626_n N_A_564_74#_c_1204_n 0.00177241f $X=6.11 $Y=1.085 $X2=0
+ $Y2=0
cc_517 N_A2_c_633_n N_A_564_74#_c_1217_n 0.00332297f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_518 N_A1_c_725_n N_VPWR_c_795_n 0.00830047f $X=6.735 $Y=1.885 $X2=0 $Y2=0
cc_519 N_A1_c_728_n N_VPWR_c_795_n 0.00787314f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_520 N_A1_c_725_n N_VPWR_c_799_n 0.00444681f $X=6.735 $Y=1.885 $X2=0 $Y2=0
cc_521 N_A1_c_728_n N_VPWR_c_800_n 0.00444681f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_522 N_A1_c_725_n N_VPWR_c_788_n 0.00429347f $X=6.735 $Y=1.885 $X2=0 $Y2=0
cc_523 N_A1_c_728_n N_VPWR_c_788_n 0.00427899f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_524 N_A1_c_725_n N_A_961_392#_c_980_n 0.00293666f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_525 N_A1_c_725_n N_A_961_392#_c_994_n 0.00233477f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_526 N_A1_c_725_n N_A_961_392#_c_998_n 0.0128308f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_527 N_A1_c_728_n N_A_961_392#_c_998_n 0.0120006f $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_528 N_A1_c_728_n N_A_961_392#_c_981_n 0.00154568f $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_529 N_A1_c_725_n N_A_1234_392#_c_1038_n 0.00542585f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_530 N_A1_c_728_n N_A_1234_392#_c_1030_n 0.00116263f $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_531 N_A1_c_729_n N_A_1234_392#_c_1030_n 4.51044e-19 $X=7.13 $Y=1.81 $X2=0
+ $Y2=0
cc_532 N_A1_c_725_n N_A_1234_392#_c_1041_n 0.0097965f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_533 N_A1_c_726_n N_A_1234_392#_c_1041_n 0.00360779f $X=6.965 $Y=1.81 $X2=0
+ $Y2=0
cc_534 N_A1_c_728_n N_A_1234_392#_c_1041_n 0.0097965f $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_535 N_A1_c_719_n N_VGND_c_1059_n 4.2194e-19 $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_536 N_A1_c_719_n N_VGND_c_1060_n 0.00356619f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_537 N_A1_c_721_n N_VGND_c_1060_n 0.00508961f $X=7.665 $Y=1.09 $X2=0 $Y2=0
cc_538 N_A1_c_719_n N_VGND_c_1067_n 0.00434272f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_539 N_A1_c_721_n N_VGND_c_1068_n 0.00434272f $X=7.665 $Y=1.09 $X2=0 $Y2=0
cc_540 N_A1_c_719_n N_VGND_c_1069_n 0.00434075f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_541 N_A1_c_721_n N_VGND_c_1069_n 0.00437635f $X=7.665 $Y=1.09 $X2=0 $Y2=0
cc_542 N_A1_c_719_n N_A_564_74#_c_1166_n 0.00668866f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_543 N_A1_c_721_n N_A_564_74#_c_1166_n 8.41862e-19 $X=7.665 $Y=1.09 $X2=0
+ $Y2=0
cc_544 N_A1_c_719_n N_A_564_74#_c_1167_n 0.0096489f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_545 N_A1_c_721_n N_A_564_74#_c_1167_n 0.0126914f $X=7.665 $Y=1.09 $X2=0 $Y2=0
cc_546 N_A1_c_722_n N_A_564_74#_c_1167_n 0.00748895f $X=7.13 $Y=1.165 $X2=0
+ $Y2=0
cc_547 N_A1_c_724_n N_A_564_74#_c_1167_n 0.0198892f $X=7.13 $Y=1.285 $X2=0 $Y2=0
cc_548 N_A1_c_719_n N_A_564_74#_c_1168_n 8.3913e-19 $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_549 N_A1_c_721_n N_A_564_74#_c_1168_n 0.00700896f $X=7.665 $Y=1.09 $X2=0
+ $Y2=0
cc_550 N_A1_c_719_n N_A_564_74#_c_1217_n 7.15802e-19 $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_551 N_A1_c_724_n N_A_564_74#_c_1217_n 0.00961222f $X=7.13 $Y=1.285 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_790_n N_X_c_887_n 7.22336e-19 $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_553 N_VPWR_c_790_n N_X_c_888_n 0.0210943f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_554 N_VPWR_c_791_n N_X_c_895_n 0.0330597f $X=1.23 $Y=2.285 $X2=0 $Y2=0
cc_555 N_VPWR_c_798_n N_X_c_895_n 0.014552f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_556 N_VPWR_c_788_n N_X_c_895_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_557 N_VPWR_M1015_d N_X_c_896_n 0.00250873f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_558 N_VPWR_c_791_n N_X_c_896_n 0.0202249f $X=1.23 $Y=2.285 $X2=0 $Y2=0
cc_559 N_VPWR_c_791_n N_X_c_897_n 0.0330597f $X=1.23 $Y=2.285 $X2=0 $Y2=0
cc_560 N_VPWR_c_792_n N_X_c_897_n 0.0146357f $X=2.085 $Y=3.33 $X2=0 $Y2=0
cc_561 N_VPWR_c_793_n N_X_c_897_n 0.0360842f $X=2.25 $Y=2.115 $X2=0 $Y2=0
cc_562 N_VPWR_c_788_n N_X_c_897_n 0.0121141f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_563 N_VPWR_c_790_n N_X_c_892_n 0.0778054f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_564 N_VPWR_c_793_n N_A_534_388#_c_962_n 0.0163153f $X=2.25 $Y=2.115 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_794_n N_A_534_388#_c_962_n 0.0116201f $X=4.36 $Y=2.79 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_796_n N_A_534_388#_c_962_n 0.0518223f $X=4.195 $Y=3.33 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_788_n N_A_534_388#_c_962_n 0.0479876f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_794_n N_A_961_392#_c_980_n 0.0182355f $X=4.36 $Y=2.79 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_795_n N_A_961_392#_c_980_n 0.00816352f $X=6.97 $Y=2.815 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_799_n N_A_961_392#_c_980_n 0.0600822f $X=6.805 $Y=3.33 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_788_n N_A_961_392#_c_980_n 0.0503539f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_572 N_VPWR_M1017_d N_A_961_392#_c_998_n 0.00427153f $X=6.81 $Y=1.96 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_795_n N_A_961_392#_c_998_n 0.0168002f $X=6.97 $Y=2.815 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_788_n N_A_961_392#_c_998_n 0.0400131f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_795_n N_A_961_392#_c_981_n 0.00681628f $X=6.97 $Y=2.815 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_800_n N_A_961_392#_c_981_n 0.0145722f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_788_n N_A_961_392#_c_981_n 0.012038f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_578 N_VPWR_M1017_d N_A_1234_392#_c_1041_n 0.00427209f $X=6.81 $Y=1.96 $X2=0
+ $Y2=0
cc_579 N_X_c_890_n N_VGND_M1019_s 0.00694709f $X=1.685 $Y=1.025 $X2=0 $Y2=0
cc_580 N_X_c_886_n N_VGND_c_1054_n 0.0126161f $X=0.685 $Y=1.225 $X2=0 $Y2=0
cc_581 N_X_c_889_n N_VGND_c_1054_n 0.0240168f $X=0.85 $Y=0.515 $X2=0 $Y2=0
cc_582 N_X_c_894_n N_VGND_c_1054_n 0.0152345f $X=0.24 $Y=1.31 $X2=0 $Y2=0
cc_583 N_X_c_889_n N_VGND_c_1055_n 0.0144922f $X=0.85 $Y=0.515 $X2=0 $Y2=0
cc_584 N_X_c_889_n N_VGND_c_1056_n 0.0165499f $X=0.85 $Y=0.515 $X2=0 $Y2=0
cc_585 N_X_c_890_n N_VGND_c_1056_n 0.0248957f $X=1.685 $Y=1.025 $X2=0 $Y2=0
cc_586 N_X_c_891_n N_VGND_c_1056_n 0.0165499f $X=1.85 $Y=0.515 $X2=0 $Y2=0
cc_587 N_X_c_891_n N_VGND_c_1057_n 0.0369264f $X=1.85 $Y=0.515 $X2=0 $Y2=0
cc_588 N_X_c_891_n N_VGND_c_1061_n 0.0145639f $X=1.85 $Y=0.515 $X2=0 $Y2=0
cc_589 N_X_c_889_n N_VGND_c_1069_n 0.0118826f $X=0.85 $Y=0.515 $X2=0 $Y2=0
cc_590 N_X_c_891_n N_VGND_c_1069_n 0.0119984f $X=1.85 $Y=0.515 $X2=0 $Y2=0
cc_591 N_A_961_392#_c_980_n N_A_1234_392#_M1010_d 0.00423003f $X=6.075 $Y=2.84
+ $X2=-0.19 $Y2=1.66
cc_592 N_A_961_392#_c_994_n N_A_1234_392#_M1010_d 0.00196975f $X=6.16 $Y=2.7
+ $X2=-0.19 $Y2=1.66
cc_593 N_A_961_392#_c_998_n N_A_1234_392#_M1010_d 0.0116068f $X=7.715 $Y=2.475
+ $X2=-0.19 $Y2=1.66
cc_594 N_A_961_392#_c_998_n N_A_1234_392#_M1018_s 0.00559058f $X=7.715 $Y=2.475
+ $X2=0 $Y2=0
cc_595 N_A_961_392#_c_998_n N_A_1234_392#_c_1031_n 0.0277488f $X=7.715 $Y=2.475
+ $X2=0 $Y2=0
cc_596 N_A_961_392#_c_991_n N_A_1234_392#_c_1031_n 0.00264697f $X=6.245 $Y=2.475
+ $X2=0 $Y2=0
cc_597 N_A_961_392#_c_982_n N_A_1234_392#_c_1030_n 0.0106894f $X=7.88 $Y=2.115
+ $X2=0 $Y2=0
cc_598 N_A_961_392#_c_998_n N_A_1234_392#_c_1041_n 0.0458302f $X=7.715 $Y=2.475
+ $X2=0 $Y2=0
cc_599 N_VGND_c_1057_n N_A_564_74#_c_1160_n 0.0346868f $X=2.405 $Y=0.515 $X2=0
+ $Y2=0
cc_600 N_VGND_c_1063_n N_A_564_74#_c_1161_n 0.0377951f $X=5.23 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_c_1069_n N_A_564_74#_c_1161_n 0.0212998f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_1057_n N_A_564_74#_c_1162_n 0.0121616f $X=2.405 $Y=0.515 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1063_n N_A_564_74#_c_1162_n 0.0235818f $X=5.23 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1069_n N_A_564_74#_c_1162_n 0.0127177f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_605 N_VGND_c_1058_n N_A_564_74#_c_1163_n 0.0100772f $X=5.395 $Y=0.525 $X2=0
+ $Y2=0
cc_606 N_VGND_c_1063_n N_A_564_74#_c_1163_n 0.065961f $X=5.23 $Y=0 $X2=0 $Y2=0
cc_607 N_VGND_c_1069_n N_A_564_74#_c_1163_n 0.0367613f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_M1000_s N_A_564_74#_c_1198_n 0.00534428f $X=5.215 $Y=0.37 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1058_n N_A_564_74#_c_1198_n 0.0203382f $X=5.395 $Y=0.525 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1069_n N_A_564_74#_c_1198_n 0.0112873f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_1058_n N_A_564_74#_c_1165_n 0.0109215f $X=5.395 $Y=0.525 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1059_n N_A_564_74#_c_1165_n 0.0105463f $X=6.395 $Y=0.52 $X2=0
+ $Y2=0
cc_613 N_VGND_c_1065_n N_A_564_74#_c_1165_n 0.0144379f $X=6.23 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_c_1069_n N_A_564_74#_c_1165_n 0.0119346f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_615 N_VGND_M1001_s N_A_564_74#_c_1208_n 0.0051536f $X=6.185 $Y=0.37 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1059_n N_A_564_74#_c_1208_n 0.0204467f $X=6.395 $Y=0.52 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1069_n N_A_564_74#_c_1208_n 0.0120866f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_618 N_VGND_c_1059_n N_A_564_74#_c_1166_n 0.0100467f $X=6.395 $Y=0.52 $X2=0
+ $Y2=0
cc_619 N_VGND_c_1060_n N_A_564_74#_c_1166_n 0.009799f $X=7.35 $Y=0.515 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1067_n N_A_564_74#_c_1166_n 0.0108951f $X=7.16 $Y=0 $X2=0 $Y2=0
cc_621 N_VGND_c_1069_n N_A_564_74#_c_1166_n 0.00900503f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_622 N_VGND_M1002_d N_A_564_74#_c_1167_n 0.00956917f $X=7.115 $Y=0.37 $X2=0
+ $Y2=0
cc_623 N_VGND_c_1060_n N_A_564_74#_c_1167_n 0.027256f $X=7.35 $Y=0.515 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1069_n N_A_564_74#_c_1167_n 0.0119957f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_625 N_VGND_c_1060_n N_A_564_74#_c_1168_n 0.0101897f $X=7.35 $Y=0.515 $X2=0
+ $Y2=0
cc_626 N_VGND_c_1068_n N_A_564_74#_c_1168_n 0.0145639f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_627 N_VGND_c_1069_n N_A_564_74#_c_1168_n 0.0119984f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_628 N_VGND_c_1063_n N_A_564_74#_c_1169_n 0.0230525f $X=5.23 $Y=0 $X2=0 $Y2=0
cc_629 N_VGND_c_1069_n N_A_564_74#_c_1169_n 0.0126179f $X=7.92 $Y=0 $X2=0 $Y2=0
