* File: sky130_fd_sc_hs__or4bb_1.pex.spice
* Created: Tue Sep  1 20:21:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__OR4BB_1%C_N 2 3 5 8 10 14 17
r32 16 17 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.52 $Y2=1.465
r33 13 16 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.29 $Y=1.465
+ $X2=0.505 $Y2=1.465
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r35 10 14 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r36 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.3 $X2=0.52
+ $Y2=1.465
r37 6 8 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.52 $Y=1.3 $X2=0.52
+ $Y2=0.645
r38 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
r39 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.955 $X2=0.505
+ $Y2=2.045
r40 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r41 1 2 126.331 $w=1.8e-07 $l=3.25e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%D_N 2 4 5 7 10 12 13 16
r53 16 18 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.215
+ $X2=1.105 $Y2=1.05
r54 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13
+ $Y=1.215 $X2=1.13 $Y2=1.215
r55 10 18 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=1.09 $Y=0.645
+ $X2=1.09 $Y2=1.05
r56 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.005 $Y=2.045
+ $X2=1.005 $Y2=2.54
r57 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.005 $Y=1.955 $X2=1.005
+ $Y2=2.045
r58 4 12 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=1.005 $Y=1.955
+ $X2=1.005 $Y2=1.72
r59 2 12 43.2981 $w=3.8e-07 $l=1.9e-07 $layer=POLY_cond $X=1.105 $Y=1.53
+ $X2=1.105 $Y2=1.72
r60 1 16 3.65891 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.105 $Y=1.24
+ $X2=1.105 $Y2=1.215
r61 1 2 42.4433 $w=3.8e-07 $l=2.9e-07 $layer=POLY_cond $X=1.105 $Y=1.24
+ $X2=1.105 $Y2=1.53
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%A_216_424# 1 2 7 9 10 12 13 20 22 26 29 31
+ 32
r65 29 31 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=1.195
+ $X2=1.695 $Y2=1.03
r66 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.74
+ $Y=1.195 $X2=1.74 $Y2=1.195
r67 24 26 5.98039 $w=5.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.305 $Y=0.615
+ $X2=1.57 $Y2=0.615
r68 22 32 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.57 $Y=1.89
+ $X2=1.57 $Y2=1.7
r69 20 32 9.97136 $w=4.18e-07 $l=2.1e-07 $layer=LI1_cond $X=1.695 $Y=1.49
+ $X2=1.695 $Y2=1.7
r70 19 29 1.23476 $w=4.18e-07 $l=4.5e-08 $layer=LI1_cond $X=1.695 $Y=1.24
+ $X2=1.695 $Y2=1.195
r71 19 20 6.85978 $w=4.18e-07 $l=2.5e-07 $layer=LI1_cond $X=1.695 $Y=1.24
+ $X2=1.695 $Y2=1.49
r72 17 26 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.57 $Y=0.88
+ $X2=1.57 $Y2=0.615
r73 17 31 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.57 $Y=0.88 $X2=1.57
+ $Y2=1.03
r74 13 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.485 $Y=2.015
+ $X2=1.57 $Y2=1.89
r75 13 15 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=1.485 $Y=2.015
+ $X2=1.34 $Y2=2.015
r76 10 30 82.0918 $w=5.74e-07 $l=7.32325e-07 $layer=POLY_cond $X=2.155 $Y=1.815
+ $X2=1.91 $Y2=1.195
r77 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.155 $Y=1.815
+ $X2=2.155 $Y2=2.39
r78 7 30 43.8845 $w=5.74e-07 $l=3.01413e-07 $layer=POLY_cond $X=2.14 $Y=1.03
+ $X2=1.91 $Y2=1.195
r79 7 9 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.14 $Y=1.03 $X2=2.14
+ $Y2=0.645
r80 2 15 600 $w=1.7e-07 $l=2.90689e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=2.12 $X2=1.34 $Y2=2.055
r81 1 24 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.165
+ $Y=0.37 $X2=1.305 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%A_27_424# 1 2 8 9 11 14 20 23 24 27 28 29 32
+ 33 36 39 42
r104 38 39 6.145 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.29
+ $X2=0.795 $Y2=2.29
r105 36 38 13.0408 $w=3.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=2.29
+ $X2=0.71 $Y2=2.29
r106 33 46 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.355
+ $X2=2.59 $Y2=1.52
r107 33 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.355
+ $X2=2.59 $Y2=1.19
r108 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.355 $X2=2.59 $Y2=1.355
r109 30 32 54.1299 $w=3.28e-07 $l=1.55e-06 $layer=LI1_cond $X=2.59 $Y=2.905
+ $X2=2.59 $Y2=1.355
r110 28 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.425 $Y=2.99
+ $X2=2.59 $Y2=2.905
r111 28 29 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.425 $Y=2.99
+ $X2=1.285 $Y2=2.99
r112 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=2.905
+ $X2=1.285 $Y2=2.99
r113 26 27 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.2 $Y=2.48
+ $X2=1.2 $Y2=2.905
r114 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=2.395
+ $X2=1.2 $Y2=2.48
r115 24 39 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.115 $Y=2.395
+ $X2=0.795 $Y2=2.395
r116 23 38 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.71 $Y=2.1 $X2=0.71
+ $Y2=2.29
r117 22 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.045
r118 22 23 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=2.1
r119 18 42 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.305 $Y=1.045
+ $X2=0.71 $Y2=1.045
r120 18 20 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.305 $Y=0.96
+ $X2=0.305 $Y2=0.645
r121 14 45 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.625 $Y=0.645
+ $X2=2.625 $Y2=1.19
r122 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.575 $Y=1.815
+ $X2=2.575 $Y2=2.39
r123 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.575 $Y=1.725
+ $X2=2.575 $Y2=1.815
r124 8 46 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.575 $Y=1.725
+ $X2=2.575 $Y2=1.52
r125 2 36 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r126 1 20 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.37 $X2=0.305 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%B 1 3 6 8 9 10 11 18
r37 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.13
+ $Y=1.515 $X2=3.13 $Y2=1.515
r38 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=2.405
+ $X2=3.13 $Y2=2.775
r39 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=2.035
+ $X2=3.13 $Y2=2.405
r40 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=1.665 $X2=3.13
+ $Y2=2.035
r41 8 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=1.515
r42 4 17 38.6549 $w=2.86e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.19 $Y=1.35
+ $X2=3.13 $Y2=1.515
r43 4 6 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.19 $Y=1.35 $X2=3.19
+ $Y2=0.645
r44 1 17 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=3.055 $Y=1.815
+ $X2=3.13 $Y2=1.515
r45 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.055 $Y=1.815
+ $X2=3.055 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%A 1 3 6 8 12
c31 6 0 2.01992e-19 $X=3.69 $Y=0.645
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.67
+ $Y=1.515 $X2=3.67 $Y2=1.515
r33 8 12 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=3.66 $Y=1.665
+ $X2=3.66 $Y2=1.515
r34 4 11 38.6549 $w=2.86e-07 $l=1.74714e-07 $layer=POLY_cond $X=3.69 $Y=1.35
+ $X2=3.67 $Y2=1.515
r35 4 6 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.69 $Y=1.35 $X2=3.69
+ $Y2=0.645
r36 1 11 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=3.595 $Y=1.815
+ $X2=3.67 $Y2=1.515
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.595 $Y=1.815
+ $X2=3.595 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%A_357_378# 1 2 3 10 12 15 23 25 29 31 34 35
+ 36 37
c88 25 0 1.25867e-19 $X=3.31 $Y=0.935
c89 10 0 3.95737e-20 $X=4.18 $Y=1.765
r90 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.465 $X2=4.21 $Y2=1.465
r91 37 38 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.475 $Y=0.935
+ $X2=3.475 $Y2=1.095
r92 34 35 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.045 $Y2=1.87
r93 32 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=1.095
+ $X2=3.475 $Y2=1.095
r94 31 42 16.3551 $w=2.76e-07 $l=4.53156e-07 $layer=LI1_cond $X=4.005 $Y=1.095
+ $X2=4.19 $Y2=1.465
r95 31 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.005 $Y=1.095
+ $X2=3.64 $Y2=1.095
r96 27 37 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0.85
+ $X2=3.475 $Y2=0.935
r97 27 29 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.475 $Y=0.85
+ $X2=3.475 $Y2=0.645
r98 26 36 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.575 $Y=0.935
+ $X2=2.325 $Y2=0.935
r99 25 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=0.935
+ $X2=3.475 $Y2=0.935
r100 25 26 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.31 $Y=0.935
+ $X2=2.575 $Y2=0.935
r101 21 36 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=0.85
+ $X2=2.325 $Y2=0.935
r102 21 23 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.41 $Y=0.85
+ $X2=2.41 $Y2=0.645
r103 19 36 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.16 $Y=1.02
+ $X2=2.325 $Y2=0.935
r104 19 35 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.16 $Y=1.02
+ $X2=2.16 $Y2=1.87
r105 13 43 38.6549 $w=2.86e-07 $l=2.03101e-07 $layer=POLY_cond $X=4.295 $Y=1.3
+ $X2=4.21 $Y2=1.465
r106 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.295 $Y=1.3
+ $X2=4.295 $Y2=0.74
r107 10 43 61.4066 $w=2.86e-07 $l=3.14643e-07 $layer=POLY_cond $X=4.18 $Y=1.765
+ $X2=4.21 $Y2=1.465
r108 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.18 $Y=1.765
+ $X2=4.18 $Y2=2.4
r109 3 34 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.785
+ $Y=1.89 $X2=1.93 $Y2=2.035
r110 2 29 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.37 $X2=3.475 $Y2=0.645
r111 1 23 182 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.37 $X2=2.41 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r46 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r48 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r49 32 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 29 32 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r54 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r58 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 20 33 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 20 30 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 18 32 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.74 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=3.33
+ $X2=3.905 $Y2=3.33
r63 17 35 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=4.56 $Y2=3.33
r64 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=3.905 $Y2=3.33
r65 13 16 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=3.905 $Y=2.115
+ $X2=3.905 $Y2=2.815
r66 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=3.245
+ $X2=3.905 $Y2=3.33
r67 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.905 $Y=3.245
+ $X2=3.905 $Y2=2.815
r68 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=3.33
r69 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=2.815
r70 2 16 600 $w=1.7e-07 $l=1.03586e-06 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=1.89 $X2=3.905 $Y2=2.815
r71 2 13 300 $w=1.7e-07 $l=3.28786e-07 $layer=licon1_PDIFF $count=2 $X=3.67
+ $Y=1.89 $X2=3.905 $Y2=2.115
r72 1 9 600 $w=1.7e-07 $l=7.88686e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.12 $X2=0.78 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%X 1 2 9 14 15 16 17 28
c23 17 0 1.15698e-19 $X=4.475 $Y=0.84
r24 21 28 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=4.53 $Y=0.945
+ $X2=4.53 $Y2=0.925
r25 17 30 8.16504 $w=3.68e-07 $l=1.53e-07 $layer=LI1_cond $X=4.53 $Y=0.977
+ $X2=4.53 $Y2=1.13
r26 17 21 0.996707 $w=3.68e-07 $l=3.2e-08 $layer=LI1_cond $X=4.53 $Y=0.977
+ $X2=4.53 $Y2=0.945
r27 17 28 1.02785 $w=3.68e-07 $l=3.3e-08 $layer=LI1_cond $X=4.53 $Y=0.892
+ $X2=4.53 $Y2=0.925
r28 16 17 11.7425 $w=3.68e-07 $l=3.77e-07 $layer=LI1_cond $X=4.53 $Y=0.515
+ $X2=4.53 $Y2=0.892
r29 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.63 $Y=1.82 $X2=4.63
+ $Y2=1.13
r30 14 15 9.3668 $w=4.73e-07 $l=1.65e-07 $layer=LI1_cond $X=4.477 $Y=1.985
+ $X2=4.477 $Y2=1.82
r31 7 14 1.813 $w=4.73e-07 $l=7.2e-08 $layer=LI1_cond $X=4.477 $Y=2.057
+ $X2=4.477 $Y2=1.985
r32 7 9 19.0869 $w=4.73e-07 $l=7.58e-07 $layer=LI1_cond $X=4.477 $Y=2.057
+ $X2=4.477 $Y2=2.815
r33 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.84 $X2=4.405 $Y2=1.985
r34 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.84 $X2=4.405 $Y2=2.815
r35 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.37
+ $Y=0.37 $X2=4.51 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_1%VGND 1 2 3 4 17 21 25 29 32 33 35 36 38 39
+ 40 53 54 57
r66 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r68 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r69 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r70 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r71 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r72 45 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r73 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.805
+ $Y2=0
r75 42 44 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.68
+ $Y2=0
r76 40 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r77 40 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r78 38 50 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.6
+ $Y2=0
r79 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.975
+ $Y2=0
r80 37 53 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.56
+ $Y2=0
r81 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=3.975
+ $Y2=0
r82 35 47 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.64
+ $Y2=0
r83 35 36 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.942
+ $Y2=0
r84 34 50 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.6
+ $Y2=0
r85 34 36 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=2.942
+ $Y2=0
r86 32 44 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.68
+ $Y2=0
r87 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.95
+ $Y2=0
r88 31 47 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.64
+ $Y2=0
r89 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=1.95
+ $Y2=0
r90 27 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=0.085
+ $X2=3.975 $Y2=0
r91 27 29 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.975 $Y=0.085
+ $X2=3.975 $Y2=0.595
r92 23 36 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.942 $Y=0.085
+ $X2=2.942 $Y2=0
r93 23 25 12.5456 $w=3.93e-07 $l=4.3e-07 $layer=LI1_cond $X=2.942 $Y=0.085
+ $X2=2.942 $Y2=0.515
r94 19 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0
r95 19 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0.515
r96 15 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0
r97 15 17 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0.57
r98 4 29 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.37 $X2=3.975 $Y2=0.595
r99 3 25 182 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.37 $X2=2.94 $Y2=0.515
r100 2 21 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.37 $X2=1.91 $Y2=0.515
r101 1 17 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.37 $X2=0.805 $Y2=0.57
.ends

