* File: sky130_fd_sc_hs__clkinv_2.pxi.spice
* Created: Thu Aug 27 20:37:05 2020
* 
x_PM_SKY130_FD_SC_HS__CLKINV_2%A N_A_M1000_g N_A_c_35_n N_A_M1002_g N_A_c_36_n
+ N_A_M1003_g N_A_c_37_n N_A_M1004_g N_A_M1001_g A A A N_A_c_34_n
+ PM_SKY130_FD_SC_HS__CLKINV_2%A
x_PM_SKY130_FD_SC_HS__CLKINV_2%Y N_Y_M1000_s N_Y_M1002_d N_Y_M1003_d N_Y_c_83_n
+ N_Y_c_84_n N_Y_c_92_n N_Y_c_85_n N_Y_c_80_n N_Y_c_86_n N_Y_c_81_n N_Y_c_105_n
+ Y PM_SKY130_FD_SC_HS__CLKINV_2%Y
x_PM_SKY130_FD_SC_HS__CLKINV_2%VPWR N_VPWR_M1002_s N_VPWR_M1004_s N_VPWR_c_130_n
+ N_VPWR_c_131_n N_VPWR_c_132_n VPWR N_VPWR_c_133_n N_VPWR_c_134_n
+ N_VPWR_c_129_n PM_SKY130_FD_SC_HS__CLKINV_2%VPWR
x_PM_SKY130_FD_SC_HS__CLKINV_2%VGND N_VGND_M1000_d N_VGND_M1001_d N_VGND_c_157_n
+ N_VGND_c_158_n N_VGND_c_159_n N_VGND_c_160_n VGND N_VGND_c_161_n
+ N_VGND_c_162_n PM_SKY130_FD_SC_HS__CLKINV_2%VGND
cc_1 VNB N_A_M1000_g 0.0644232f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_2 VNB N_A_M1001_g 0.0581471f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.61
cc_3 VNB A 0.0183006f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_A_c_34_n 0.0669284f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.557
cc_5 VNB N_Y_c_80_n 0.0153843f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_6 VNB N_Y_c_81_n 0.0174246f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.557
cc_7 VNB Y 0.0240108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_VPWR_c_129_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.557
cc_9 VNB N_VGND_c_157_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_10 VNB N_VGND_c_158_n 0.0338694f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_11 VNB N_VGND_c_159_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.765
cc_12 VNB N_VGND_c_160_n 0.0321896f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_13 VNB N_VGND_c_161_n 0.0287859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_162_n 0.143782f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_15 VPB N_A_c_35_n 0.0208611f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_16 VPB N_A_c_36_n 0.0155104f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_17 VPB N_A_c_37_n 0.0163707f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_18 VPB A 0.0143109f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_19 VPB N_A_c_34_n 0.0351528f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.557
cc_20 VPB N_Y_c_83_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_21 VPB N_Y_c_84_n 0.0353617f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_22 VPB N_Y_c_85_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_23 VPB N_Y_c_86_n 0.00714919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_24 VPB Y 0.01299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_25 VPB N_VPWR_c_130_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_26 VPB N_VPWR_c_131_n 0.0108116f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_27 VPB N_VPWR_c_132_n 0.0370539f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.61
cc_28 VPB N_VPWR_c_133_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_29 VPB N_VPWR_c_134_n 0.0234893f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.557
cc_30 VPB N_VPWR_c_129_n 0.0580979f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.557
cc_31 N_A_c_35_n N_Y_c_83_n 4.27055e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_32 A N_Y_c_83_n 0.0260502f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_33 N_A_c_35_n N_Y_c_84_n 0.0104891f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_34 N_A_c_36_n N_Y_c_84_n 6.45594e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_35 N_A_c_35_n N_Y_c_92_n 0.0120074f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_36 N_A_c_36_n N_Y_c_92_n 0.0120074f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_37 A N_Y_c_92_n 0.0393875f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_38 N_A_c_34_n N_Y_c_92_n 0.00131635f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_39 N_A_c_35_n N_Y_c_85_n 6.45594e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_40 N_A_c_36_n N_Y_c_85_n 0.0103431f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_41 N_A_c_37_n N_Y_c_85_n 0.01498f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_42 N_A_M1001_g N_Y_c_80_n 0.0222952f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_43 N_A_c_37_n N_Y_c_86_n 0.0173803f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_44 N_A_M1000_g N_Y_c_81_n 0.0223806f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_45 N_A_M1001_g N_Y_c_81_n 0.0144176f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_46 A N_Y_c_81_n 0.0596487f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_47 N_A_c_34_n N_Y_c_81_n 0.014563f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_48 N_A_c_36_n N_Y_c_105_n 4.27055e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_49 N_A_c_37_n N_Y_c_105_n 9.50925e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_50 A N_Y_c_105_n 0.0217109f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_51 N_A_c_34_n N_Y_c_105_n 0.00143147f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_52 N_A_c_37_n Y 0.00697061f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_53 N_A_M1001_g Y 0.0190699f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_54 A Y 0.0265979f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_55 N_A_c_35_n N_VPWR_c_130_n 0.00486623f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_56 N_A_c_36_n N_VPWR_c_130_n 0.00486623f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A_c_37_n N_VPWR_c_132_n 0.00714506f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_58 N_A_c_36_n N_VPWR_c_133_n 0.00445602f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_59 N_A_c_37_n N_VPWR_c_133_n 0.00445602f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_60 N_A_c_35_n N_VPWR_c_134_n 0.00445602f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A_c_35_n N_VPWR_c_129_n 0.008611f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A_c_36_n N_VPWR_c_129_n 0.00857589f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_63 N_A_c_37_n N_VPWR_c_129_n 0.008611f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_VGND_c_158_n 0.0187336f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_65 A N_VGND_c_158_n 0.013195f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_66 N_A_M1001_g N_VGND_c_160_n 0.0184421f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_VGND_c_161_n 0.00462012f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_68 N_A_M1001_g N_VGND_c_161_n 0.00462012f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_69 N_A_M1000_g N_VGND_c_162_n 0.00450456f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_70 N_A_M1001_g N_VGND_c_162_n 0.00450456f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_71 N_Y_c_92_n N_VPWR_M1002_s 0.00408911f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_72 N_Y_c_86_n N_VPWR_M1004_s 0.00477129f $X=1.565 $Y=2.035 $X2=0 $Y2=0
cc_73 Y N_VPWR_M1004_s 0.00194528f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_74 N_Y_c_84_n N_VPWR_c_130_n 0.0449718f $X=0.285 $Y=2.815 $X2=0 $Y2=0
cc_75 N_Y_c_92_n N_VPWR_c_130_n 0.0136682f $X=1.02 $Y=2.035 $X2=0 $Y2=0
cc_76 N_Y_c_85_n N_VPWR_c_130_n 0.0449718f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_77 N_Y_c_85_n N_VPWR_c_132_n 0.0462948f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_78 N_Y_c_86_n N_VPWR_c_132_n 0.0218009f $X=1.565 $Y=2.035 $X2=0 $Y2=0
cc_79 N_Y_c_85_n N_VPWR_c_133_n 0.014552f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_80 N_Y_c_84_n N_VPWR_c_134_n 0.0145938f $X=0.285 $Y=2.815 $X2=0 $Y2=0
cc_81 N_Y_c_84_n N_VPWR_c_129_n 0.0120466f $X=0.285 $Y=2.815 $X2=0 $Y2=0
cc_82 N_Y_c_85_n N_VPWR_c_129_n 0.0119791f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_83 N_Y_c_81_n N_VGND_c_158_n 0.0132912f $X=1.305 $Y=0.845 $X2=0 $Y2=0
cc_84 N_Y_c_80_n N_VGND_c_160_n 0.0288308f $X=1.565 $Y=1.095 $X2=0 $Y2=0
cc_85 N_Y_c_81_n N_VGND_c_160_n 0.0132912f $X=1.305 $Y=0.845 $X2=0 $Y2=0
cc_86 N_Y_c_81_n N_VGND_c_161_n 0.0175309f $X=1.305 $Y=0.845 $X2=0 $Y2=0
cc_87 N_Y_c_81_n N_VGND_c_162_n 0.0228888f $X=1.305 $Y=0.845 $X2=0 $Y2=0
