* NGSPICE file created from sky130_fd_sc_hs__tapmet1_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__tapmet1_2 VGND VPB VPWR
.ends

