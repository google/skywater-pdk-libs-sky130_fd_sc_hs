* File: sky130_fd_sc_hs__o41ai_4.pxi.spice
* Created: Tue Sep  1 20:19:41 2020
* 
x_PM_SKY130_FD_SC_HS__O41AI_4%B1 N_B1_c_149_n N_B1_M1017_g N_B1_c_156_n
+ N_B1_M1015_g N_B1_c_150_n N_B1_M1022_g N_B1_c_157_n N_B1_M1026_g N_B1_c_151_n
+ N_B1_M1030_g N_B1_c_152_n N_B1_c_153_n N_B1_c_154_n N_B1_M1031_g B1 B1
+ N_B1_c_155_n PM_SKY130_FD_SC_HS__O41AI_4%B1
x_PM_SKY130_FD_SC_HS__O41AI_4%A4 N_A4_c_223_n N_A4_M1000_g N_A4_c_216_n
+ N_A4_M1002_g N_A4_c_224_n N_A4_M1004_g N_A4_c_225_n N_A4_M1029_g N_A4_c_217_n
+ N_A4_M1012_g N_A4_c_226_n N_A4_M1035_g N_A4_c_218_n N_A4_M1024_g N_A4_c_219_n
+ N_A4_c_220_n N_A4_c_221_n N_A4_M1027_g A4 A4 N_A4_c_222_n
+ PM_SKY130_FD_SC_HS__O41AI_4%A4
x_PM_SKY130_FD_SC_HS__O41AI_4%A3 N_A3_c_312_n N_A3_M1001_g N_A3_c_304_n
+ N_A3_c_305_n N_A3_c_306_n N_A3_M1003_g N_A3_c_315_n N_A3_M1006_g N_A3_c_316_n
+ N_A3_M1007_g N_A3_c_307_n N_A3_M1032_g N_A3_c_317_n N_A3_M1014_g N_A3_c_308_n
+ N_A3_M1036_g N_A3_c_309_n N_A3_M1037_g A3 A3 A3 A3 N_A3_c_311_n
+ PM_SKY130_FD_SC_HS__O41AI_4%A3
x_PM_SKY130_FD_SC_HS__O41AI_4%A2 N_A2_c_408_n N_A2_M1005_g N_A2_c_414_n
+ N_A2_M1009_g N_A2_c_409_n N_A2_M1023_g N_A2_c_415_n N_A2_M1010_g N_A2_c_410_n
+ N_A2_M1025_g N_A2_c_416_n N_A2_M1013_g N_A2_c_411_n N_A2_M1028_g N_A2_c_417_n
+ N_A2_M1016_g A2 A2 A2 A2 N_A2_c_413_n PM_SKY130_FD_SC_HS__O41AI_4%A2
x_PM_SKY130_FD_SC_HS__O41AI_4%A1 N_A1_c_509_n N_A1_M1018_g N_A1_c_503_n
+ N_A1_M1008_g N_A1_c_510_n N_A1_M1019_g N_A1_c_504_n N_A1_M1011_g N_A1_c_511_n
+ N_A1_M1020_g N_A1_c_505_n N_A1_M1033_g N_A1_c_512_n N_A1_M1021_g N_A1_c_506_n
+ N_A1_M1034_g A1 A1 A1 A1 N_A1_c_508_n PM_SKY130_FD_SC_HS__O41AI_4%A1
x_PM_SKY130_FD_SC_HS__O41AI_4%VPWR N_VPWR_M1015_d N_VPWR_M1026_d N_VPWR_M1018_s
+ N_VPWR_M1020_s N_VPWR_c_582_n N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n
+ N_VPWR_c_586_n VPWR N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n
+ N_VPWR_c_590_n N_VPWR_c_581_n N_VPWR_c_592_n N_VPWR_c_593_n N_VPWR_c_594_n
+ PM_SKY130_FD_SC_HS__O41AI_4%VPWR
x_PM_SKY130_FD_SC_HS__O41AI_4%Y N_Y_M1017_s N_Y_M1030_s N_Y_M1015_s N_Y_M1000_d
+ N_Y_M1029_d N_Y_c_689_n N_Y_c_698_n N_Y_c_690_n N_Y_c_691_n N_Y_c_708_n
+ N_Y_c_688_n N_Y_c_693_n N_Y_c_745_p N_Y_c_694_n N_Y_c_748_p N_Y_c_715_n
+ N_Y_c_695_n N_Y_c_726_n Y Y N_Y_c_728_n PM_SKY130_FD_SC_HS__O41AI_4%Y
x_PM_SKY130_FD_SC_HS__O41AI_4%A_339_368# N_A_339_368#_M1000_s
+ N_A_339_368#_M1004_s N_A_339_368#_M1035_s N_A_339_368#_M1006_d
+ N_A_339_368#_M1014_d N_A_339_368#_c_760_n N_A_339_368#_c_761_n
+ N_A_339_368#_c_762_n N_A_339_368#_c_775_n N_A_339_368#_c_763_n
+ N_A_339_368#_c_764_n N_A_339_368#_c_765_n N_A_339_368#_c_785_n
+ N_A_339_368#_c_766_n N_A_339_368#_c_767_n N_A_339_368#_c_768_n
+ N_A_339_368#_c_769_n N_A_339_368#_c_770_n
+ PM_SKY130_FD_SC_HS__O41AI_4%A_339_368#
x_PM_SKY130_FD_SC_HS__O41AI_4%A_788_368# N_A_788_368#_M1001_s
+ N_A_788_368#_M1007_s N_A_788_368#_M1009_d N_A_788_368#_M1013_d
+ N_A_788_368#_c_871_n N_A_788_368#_c_845_n N_A_788_368#_c_841_n
+ N_A_788_368#_c_875_n N_A_788_368#_c_842_n N_A_788_368#_c_882_p
+ N_A_788_368#_c_843_n N_A_788_368#_c_885_p N_A_788_368#_c_856_n
+ N_A_788_368#_c_844_n PM_SKY130_FD_SC_HS__O41AI_4%A_788_368#
x_PM_SKY130_FD_SC_HS__O41AI_4%A_1191_368# N_A_1191_368#_M1009_s
+ N_A_1191_368#_M1010_s N_A_1191_368#_M1016_s N_A_1191_368#_M1019_d
+ N_A_1191_368#_M1021_d N_A_1191_368#_c_888_n N_A_1191_368#_c_889_n
+ N_A_1191_368#_c_890_n N_A_1191_368#_c_906_n N_A_1191_368#_c_891_n
+ N_A_1191_368#_c_912_n N_A_1191_368#_c_892_n N_A_1191_368#_c_893_n
+ N_A_1191_368#_c_894_n N_A_1191_368#_c_895_n N_A_1191_368#_c_896_n
+ N_A_1191_368#_c_897_n N_A_1191_368#_c_898_n
+ PM_SKY130_FD_SC_HS__O41AI_4%A_1191_368#
x_PM_SKY130_FD_SC_HS__O41AI_4%A_27_74# N_A_27_74#_M1017_d N_A_27_74#_M1022_d
+ N_A_27_74#_M1031_d N_A_27_74#_M1012_s N_A_27_74#_M1027_s N_A_27_74#_M1032_s
+ N_A_27_74#_M1037_s N_A_27_74#_M1023_d N_A_27_74#_M1028_d N_A_27_74#_M1011_d
+ N_A_27_74#_M1034_d N_A_27_74#_c_970_n N_A_27_74#_c_971_n N_A_27_74#_c_972_n
+ N_A_27_74#_c_973_n N_A_27_74#_c_1001_n N_A_27_74#_c_1002_n N_A_27_74#_c_1006_n
+ N_A_27_74#_c_974_n N_A_27_74#_c_975_n N_A_27_74#_c_976_n N_A_27_74#_c_1017_n
+ N_A_27_74#_c_977_n N_A_27_74#_c_978_n N_A_27_74#_c_1033_n N_A_27_74#_c_979_n
+ N_A_27_74#_c_1040_n N_A_27_74#_c_980_n N_A_27_74#_c_1053_n N_A_27_74#_c_981_n
+ N_A_27_74#_c_1059_n N_A_27_74#_c_982_n N_A_27_74#_c_1069_n N_A_27_74#_c_983_n
+ N_A_27_74#_c_1077_n N_A_27_74#_c_984_n N_A_27_74#_c_985_n N_A_27_74#_c_986_n
+ N_A_27_74#_c_1022_n N_A_27_74#_c_1024_n N_A_27_74#_c_1047_n
+ N_A_27_74#_c_1050_n N_A_27_74#_c_1065_n N_A_27_74#_c_1067_n
+ N_A_27_74#_c_1083_n PM_SKY130_FD_SC_HS__O41AI_4%A_27_74#
x_PM_SKY130_FD_SC_HS__O41AI_4%VGND N_VGND_M1002_d N_VGND_M1024_d N_VGND_M1003_d
+ N_VGND_M1036_d N_VGND_M1005_s N_VGND_M1025_s N_VGND_M1008_s N_VGND_M1033_s
+ N_VGND_c_1160_n N_VGND_c_1161_n N_VGND_c_1162_n N_VGND_c_1163_n
+ N_VGND_c_1164_n N_VGND_c_1165_n N_VGND_c_1166_n N_VGND_c_1167_n
+ N_VGND_c_1168_n N_VGND_c_1169_n N_VGND_c_1170_n VGND N_VGND_c_1171_n
+ N_VGND_c_1172_n N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n
+ N_VGND_c_1176_n N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n
+ N_VGND_c_1180_n N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n
+ PM_SKY130_FD_SC_HS__O41AI_4%VGND
cc_1 VNB N_B1_c_149_n 0.0185832f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_2 VNB N_B1_c_150_n 0.0143157f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.185
cc_3 VNB N_B1_c_151_n 0.0149371f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.185
cc_4 VNB N_B1_c_152_n 0.0298945f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.26
cc_5 VNB N_B1_c_153_n 0.111235f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.26
cc_6 VNB N_B1_c_154_n 0.0152736f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.185
cc_7 VNB N_B1_c_155_n 0.0259935f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.385
cc_8 VNB N_A4_c_216_n 0.0173669f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_9 VNB N_A4_c_217_n 0.0173529f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.185
cc_10 VNB N_A4_c_218_n 0.0151591f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_11 VNB N_A4_c_219_n 0.0185585f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_A4_c_220_n 0.120189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A4_c_221_n 0.0151037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A4_c_222_n 0.0115136f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_15 VNB N_A3_c_304_n 0.0119481f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_16 VNB N_A3_c_305_n 0.00654076f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_17 VNB N_A3_c_306_n 0.0178826f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB N_A3_c_307_n 0.0168239f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_19 VNB N_A3_c_308_n 0.0173859f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_A3_c_309_n 0.0171629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A3 0.0173798f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.475
cc_22 VNB N_A3_c_311_n 0.113713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_c_408_n 0.0180414f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_24 VNB N_A2_c_409_n 0.0168231f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.185
cc_25 VNB N_A2_c_410_n 0.0165146f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.185
cc_26 VNB N_A2_c_411_n 0.0179931f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_27 VNB A2 0.0177499f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_28 VNB N_A2_c_413_n 0.11479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_c_503_n 0.0181973f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_30 VNB N_A1_c_504_n 0.0175147f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.765
cc_31 VNB N_A1_c_505_n 0.0173888f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.26
cc_32 VNB N_A1_c_506_n 0.0228112f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_33 VNB A1 0.0307917f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_34 VNB N_A1_c_508_n 0.12313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_581_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_688_n 0.00830153f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.385
cc_37 VNB N_A_27_74#_c_970_n 0.0226322f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_38 VNB N_A_27_74#_c_971_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_972_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.365
cc_40 VNB N_A_27_74#_c_973_n 0.00502562f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_41 VNB N_A_27_74#_c_974_n 0.0028074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_975_n 6.81442e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_976_n 0.00753795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_74#_c_977_n 0.00240128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_74#_c_978_n 0.00140577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_74#_c_979_n 0.00206561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_980_n 0.00206561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_981_n 0.00178829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_74#_c_982_n 0.00253253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_74#_c_983_n 0.0024006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_27_74#_c_984_n 0.0075085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_74#_c_985_n 0.0203664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_27_74#_c_986_n 0.00202117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1160_n 0.00933987f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.385
cc_55 VNB N_VGND_c_1161_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.475
cc_56 VNB N_VGND_c_1162_n 0.00578139f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.385
cc_57 VNB N_VGND_c_1163_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.185
cc_58 VNB N_VGND_c_1164_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.365
cc_59 VNB N_VGND_c_1165_n 0.00485164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1166_n 0.00498382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1167_n 0.00528272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1168_n 0.00571618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1169_n 0.0189539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1170_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1171_n 0.0809332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1172_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1173_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1174_n 0.018048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1175_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1176_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1177_n 0.507588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1178_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1179_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1180_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1181_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1182_n 0.00617178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1183_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VPB N_B1_c_156_n 0.0194239f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_79 VPB N_B1_c_157_n 0.0181146f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.765
cc_80 VPB N_B1_c_153_n 0.0180757f $X=-0.19 $Y=1.66 $X2=1.43 $Y2=1.26
cc_81 VPB N_A4_c_223_n 0.0170303f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_82 VPB N_A4_c_224_n 0.0141098f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.185
cc_83 VPB N_A4_c_225_n 0.0141098f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.765
cc_84 VPB N_A4_c_226_n 0.0148744f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.26
cc_85 VPB N_A4_c_220_n 0.0485666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A3_c_312_n 0.0153478f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_87 VPB N_A3_c_304_n 0.0133997f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_88 VPB N_A3_c_305_n 0.00590087f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_89 VPB N_A3_c_315_n 0.014812f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_90 VPB N_A3_c_316_n 0.0141056f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.4
cc_91 VPB N_A3_c_317_n 0.0172095f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.185
cc_92 VPB N_A3_c_311_n 0.0349113f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A2_c_414_n 0.0172095f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_94 VPB N_A2_c_415_n 0.0141056f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.765
cc_95 VPB N_A2_c_416_n 0.0141056f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.26
cc_96 VPB N_A2_c_417_n 0.0144441f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_97 VPB N_A2_c_413_n 0.0275577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A1_c_509_n 0.0149969f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_99 VPB N_A1_c_510_n 0.0152448f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.185
cc_100 VPB N_A1_c_511_n 0.0152448f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.185
cc_101 VPB N_A1_c_512_n 0.0185559f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=0.74
cc_102 VPB N_A1_c_508_n 0.0278339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_582_n 0.0120106f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.185
cc_104 VPB N_VPWR_c_583_n 0.0556112f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_105 VPB N_VPWR_c_584_n 0.0141288f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_106 VPB N_VPWR_c_585_n 0.00575879f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.475
cc_107 VPB N_VPWR_c_586_n 0.00575879f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.475
cc_108 VPB N_VPWR_c_587_n 0.0183788f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.385
cc_109 VPB N_VPWR_c_588_n 0.155087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_589_n 0.0185924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_590_n 0.0177062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_581_n 0.111616f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_592_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_593_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_594_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_Y_c_689_n 0.00326535f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.185
cc_117 VPB N_Y_c_690_n 0.0059192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_Y_c_691_n 0.00432492f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.475
cc_119 VPB N_Y_c_688_n 0.00201193f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.385
cc_120 VPB N_Y_c_693_n 0.00297633f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.475
cc_121 VPB N_Y_c_694_n 5.66347e-19 $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.475
cc_122 VPB N_Y_c_695_n 0.0101507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_339_368#_c_760_n 0.00766789f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.185
cc_124 VPB N_A_339_368#_c_761_n 0.00226419f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=0.74
cc_125 VPB N_A_339_368#_c_762_n 0.00424176f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_126 VPB N_A_339_368#_c_763_n 0.00226419f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.385
cc_127 VPB N_A_339_368#_c_764_n 0.00294354f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.475
cc_128 VPB N_A_339_368#_c_765_n 0.0030167f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.475
cc_129 VPB N_A_339_368#_c_766_n 0.00644841f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_130 VPB N_A_339_368#_c_767_n 0.00763926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_339_368#_c_768_n 0.00203831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_339_368#_c_769_n 0.00211111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_339_368#_c_770_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_788_368#_c_841_n 9.52341e-19 $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.185
cc_135 VPB N_A_788_368#_c_842_n 0.0188562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_788_368#_c_843_n 0.0053512f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.475
cc_137 VPB N_A_788_368#_c_844_n 0.00186725f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_138 VPB N_A_1191_368#_c_888_n 0.00754475f $X=-0.19 $Y=1.66 $X2=1.855
+ $Y2=1.185
cc_139 VPB N_A_1191_368#_c_889_n 0.00213916f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=0.74
cc_140 VPB N_A_1191_368#_c_890_n 0.00444759f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_141 VPB N_A_1191_368#_c_891_n 0.00506057f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.385
cc_142 VPB N_A_1191_368#_c_892_n 0.00443091f $X=-0.19 $Y=1.66 $X2=1.055
+ $Y2=1.475
cc_143 VPB N_A_1191_368#_c_893_n 0.00234762f $X=-0.19 $Y=1.66 $X2=1.355
+ $Y2=1.185
cc_144 VPB N_A_1191_368#_c_894_n 0.00248717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1191_368#_c_895_n 0.0131052f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.365
cc_146 VPB N_A_1191_368#_c_896_n 0.0441891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_1191_368#_c_897_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1191_368#_c_898_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 N_B1_c_154_n N_A4_c_216_n 0.0177689f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_150 N_B1_c_152_n N_A4_c_220_n 0.00932861f $X=1.78 $Y=1.26 $X2=0 $Y2=0
cc_151 N_B1_c_154_n N_A4_c_222_n 0.00137652f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_152 N_B1_c_156_n N_VPWR_c_583_n 0.0178484f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_153 N_B1_c_157_n N_VPWR_c_583_n 6.08597e-19 $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_154 N_B1_c_153_n N_VPWR_c_583_n 0.00677955f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_155 N_B1_c_155_n N_VPWR_c_583_n 0.0191836f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_156 N_B1_c_156_n N_VPWR_c_584_n 5.26157e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_157 N_B1_c_157_n N_VPWR_c_584_n 0.0181585f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B1_c_156_n N_VPWR_c_587_n 0.00413917f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B1_c_157_n N_VPWR_c_587_n 0.00413917f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_160 N_B1_c_156_n N_VPWR_c_581_n 0.00818606f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_161 N_B1_c_157_n N_VPWR_c_581_n 0.00818606f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B1_c_156_n N_Y_c_689_n 0.0065528f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B1_c_157_n N_Y_c_689_n 0.0065528f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B1_c_150_n N_Y_c_698_n 0.00955428f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_165 N_B1_c_151_n N_Y_c_698_n 0.015868f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_166 N_B1_c_153_n N_Y_c_698_n 0.00191032f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_167 N_B1_c_155_n N_Y_c_698_n 0.0224794f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_168 N_B1_c_157_n N_Y_c_690_n 0.0126105f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B1_c_153_n N_Y_c_690_n 0.0159661f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_170 N_B1_c_155_n N_Y_c_690_n 0.0144526f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_171 N_B1_c_156_n N_Y_c_691_n 0.00235826f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_172 N_B1_c_153_n N_Y_c_691_n 0.00646827f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_173 N_B1_c_155_n N_Y_c_691_n 0.0280525f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_174 N_B1_c_154_n N_Y_c_708_n 0.0054601f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_175 N_B1_c_151_n N_Y_c_688_n 0.00255143f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_176 N_B1_c_152_n N_Y_c_688_n 0.0205092f $X=1.78 $Y=1.26 $X2=0 $Y2=0
cc_177 N_B1_c_153_n N_Y_c_688_n 0.00684117f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_178 N_B1_c_154_n N_Y_c_688_n 0.0048483f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_179 N_B1_c_155_n N_Y_c_688_n 0.0181698f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_180 N_B1_c_152_n N_Y_c_693_n 0.00411697f $X=1.78 $Y=1.26 $X2=0 $Y2=0
cc_181 N_B1_c_153_n N_Y_c_715_n 7.43006e-19 $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_182 N_B1_c_155_n N_Y_c_715_n 0.0140705f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_183 N_B1_c_157_n N_A_339_368#_c_760_n 0.00184524f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_B1_c_157_n N_A_339_368#_c_762_n 5.94256e-19 $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_B1_c_149_n N_A_27_74#_c_970_n 0.00796844f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_186 N_B1_c_150_n N_A_27_74#_c_970_n 5.73078e-19 $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_187 N_B1_c_153_n N_A_27_74#_c_970_n 0.00205263f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_188 N_B1_c_155_n N_A_27_74#_c_970_n 0.0251377f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_189 N_B1_c_149_n N_A_27_74#_c_971_n 0.0100711f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_190 N_B1_c_150_n N_A_27_74#_c_971_n 0.00789822f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_191 N_B1_c_149_n N_A_27_74#_c_972_n 0.00282152f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_192 N_B1_c_151_n N_A_27_74#_c_973_n 0.00829147f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_193 N_B1_c_154_n N_A_27_74#_c_973_n 0.0137299f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_194 N_B1_c_149_n N_A_27_74#_c_986_n 6.04287e-19 $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_195 N_B1_c_150_n N_A_27_74#_c_986_n 0.00642184f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_196 N_B1_c_151_n N_A_27_74#_c_986_n 0.00684618f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_197 N_B1_c_154_n N_A_27_74#_c_986_n 6.66855e-19 $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_198 N_B1_c_149_n N_VGND_c_1171_n 0.00278247f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_199 N_B1_c_150_n N_VGND_c_1171_n 0.00279469f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_200 N_B1_c_151_n N_VGND_c_1171_n 0.00279469f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_201 N_B1_c_154_n N_VGND_c_1171_n 0.00278271f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_202 N_B1_c_149_n N_VGND_c_1177_n 0.00357084f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_203 N_B1_c_150_n N_VGND_c_1177_n 0.00352518f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_204 N_B1_c_151_n N_VGND_c_1177_n 0.00353176f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_205 N_B1_c_154_n N_VGND_c_1177_n 0.00354798f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_206 N_A4_c_226_n N_A3_c_312_n 0.0114755f $X=3.415 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_207 N_A4_c_219_n N_A3_c_305_n 0.0142465f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_208 N_A4_c_220_n N_A3_c_305_n 0.0117084f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_209 N_A4_c_221_n N_A3_c_306_n 0.00804366f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_210 N_A4_c_219_n N_A3_c_311_n 0.00804366f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_211 N_A4_c_223_n N_VPWR_c_584_n 8.67856e-19 $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A4_c_223_n N_VPWR_c_588_n 0.00278271f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A4_c_224_n N_VPWR_c_588_n 0.00278271f $X=2.515 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A4_c_225_n N_VPWR_c_588_n 0.00278271f $X=2.965 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A4_c_226_n N_VPWR_c_588_n 0.00278271f $X=3.415 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A4_c_223_n N_VPWR_c_581_n 0.00358624f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A4_c_224_n N_VPWR_c_581_n 0.00353823f $X=2.515 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A4_c_225_n N_VPWR_c_581_n 0.00353823f $X=2.965 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A4_c_226_n N_VPWR_c_581_n 0.00353907f $X=3.415 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A4_c_216_n N_Y_c_688_n 5.71389e-19 $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_221 N_A4_c_220_n N_Y_c_688_n 0.00868138f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_222 N_A4_c_222_n N_Y_c_688_n 0.0248693f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_223 N_A4_c_223_n N_Y_c_693_n 0.01221f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A4_c_220_n N_Y_c_693_n 0.00571116f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_225 N_A4_c_222_n N_Y_c_693_n 0.00796928f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_226 N_A4_c_226_n N_Y_c_694_n 9.86303e-19 $X=3.415 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A4_c_220_n N_Y_c_694_n 0.0191305f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_228 N_A4_c_222_n N_Y_c_694_n 0.00885397f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_229 N_A4_c_220_n N_Y_c_726_n 0.0121675f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_230 N_A4_c_222_n N_Y_c_726_n 0.0225374f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_231 N_A4_c_224_n N_Y_c_728_n 0.0184885f $X=2.515 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A4_c_225_n N_Y_c_728_n 0.0183458f $X=2.965 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A4_c_220_n N_Y_c_728_n 0.0181766f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_234 N_A4_c_222_n N_Y_c_728_n 0.0478219f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_235 N_A4_c_223_n N_A_339_368#_c_761_n 0.0141328f $X=2.065 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A4_c_224_n N_A_339_368#_c_761_n 0.0132631f $X=2.515 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A4_c_220_n N_A_339_368#_c_775_n 7.81626e-19 $X=3.615 $Y=1.26 $X2=0
+ $Y2=0
cc_238 N_A4_c_225_n N_A_339_368#_c_763_n 0.0132631f $X=2.965 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A4_c_226_n N_A_339_368#_c_763_n 0.0132287f $X=3.415 $Y=1.765 $X2=0
+ $Y2=0
cc_240 N_A4_c_226_n N_A_339_368#_c_764_n 7.74287e-19 $X=3.415 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A4_c_220_n N_A_339_368#_c_764_n 0.00152953f $X=3.615 $Y=1.26 $X2=0
+ $Y2=0
cc_242 N_A4_c_216_n N_A_27_74#_c_973_n 0.00353966f $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_243 N_A4_c_216_n N_A_27_74#_c_1001_n 0.0124539f $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_244 N_A4_c_216_n N_A_27_74#_c_1002_n 0.00979933f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_245 N_A4_c_217_n N_A_27_74#_c_1002_n 0.0111145f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_246 N_A4_c_220_n N_A_27_74#_c_1002_n 0.00275601f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_247 N_A4_c_222_n N_A_27_74#_c_1002_n 0.0612456f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_248 N_A4_c_216_n N_A_27_74#_c_1006_n 7.32094e-19 $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_249 N_A4_c_220_n N_A_27_74#_c_1006_n 0.00298138f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_250 N_A4_c_222_n N_A_27_74#_c_1006_n 0.0199556f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_251 N_A4_c_217_n N_A_27_74#_c_974_n 2.68164e-19 $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_252 N_A4_c_218_n N_A_27_74#_c_974_n 0.00604445f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_253 N_A4_c_217_n N_A_27_74#_c_975_n 0.0032036f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_254 N_A4_c_218_n N_A_27_74#_c_975_n 0.00281435f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_255 N_A4_c_220_n N_A_27_74#_c_975_n 0.00726061f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_256 N_A4_c_222_n N_A_27_74#_c_975_n 0.00900371f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_257 N_A4_c_219_n N_A_27_74#_c_976_n 0.018043f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_258 N_A4_c_220_n N_A_27_74#_c_976_n 0.0105089f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_259 N_A4_c_220_n N_A_27_74#_c_1017_n 0.0138097f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_260 N_A4_c_222_n N_A_27_74#_c_1017_n 0.0143906f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_261 N_A4_c_221_n N_A_27_74#_c_977_n 0.00574886f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_262 N_A4_c_219_n N_A_27_74#_c_978_n 0.00388347f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_263 N_A4_c_221_n N_A_27_74#_c_978_n 0.00267912f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_264 N_A4_c_218_n N_A_27_74#_c_1022_n 0.00184154f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_265 N_A4_c_220_n N_A_27_74#_c_1022_n 0.00369173f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_266 N_A4_c_221_n N_A_27_74#_c_1024_n 0.0017646f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_267 N_A4_c_218_n N_VGND_c_1160_n 0.00313396f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_268 N_A4_c_219_n N_VGND_c_1160_n 0.00230361f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_269 N_A4_c_221_n N_VGND_c_1160_n 0.00313962f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_270 N_A4_c_221_n N_VGND_c_1161_n 0.00434272f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_271 N_A4_c_217_n N_VGND_c_1169_n 0.00461464f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_272 N_A4_c_218_n N_VGND_c_1169_n 0.00422942f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_273 N_A4_c_216_n N_VGND_c_1171_n 0.00789845f $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_274 N_A4_c_217_n N_VGND_c_1171_n 0.00590535f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_275 N_A4_c_216_n N_VGND_c_1177_n 0.00447853f $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_276 N_A4_c_217_n N_VGND_c_1177_n 0.00465356f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A4_c_218_n N_VGND_c_1177_n 0.00783843f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_278 N_A4_c_221_n N_VGND_c_1177_n 0.00820382f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_279 N_A3_c_309_n N_A2_c_408_n 0.00936575f $X=5.83 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_280 A3 N_A2_c_408_n 0.0044767f $X=5.915 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_281 A3 A2 0.0247108f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_282 N_A3_c_311_n A2 2.21735e-19 $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_283 N_A3_c_311_n N_A2_c_413_n 0.0132359f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_284 N_A3_c_312_n N_VPWR_c_588_n 0.00278257f $X=3.865 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A3_c_315_n N_VPWR_c_588_n 0.00278257f $X=4.415 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A3_c_316_n N_VPWR_c_588_n 0.00278257f $X=4.865 $Y=1.765 $X2=0 $Y2=0
cc_287 N_A3_c_317_n N_VPWR_c_588_n 0.00278257f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A3_c_312_n N_VPWR_c_581_n 0.00354785f $X=3.865 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A3_c_315_n N_VPWR_c_581_n 0.00354701f $X=4.415 $Y=1.765 $X2=0 $Y2=0
cc_290 N_A3_c_316_n N_VPWR_c_581_n 0.00353822f $X=4.865 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A3_c_317_n N_VPWR_c_581_n 0.00358623f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A3_c_312_n N_A_339_368#_c_764_n 0.0138585f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A3_c_305_n N_A_339_368#_c_764_n 4.19419e-19 $X=3.955 $Y=1.65 $X2=0
+ $Y2=0
cc_294 N_A3_c_315_n N_A_339_368#_c_764_n 7.56633e-19 $X=4.415 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A3_c_312_n N_A_339_368#_c_765_n 0.0113536f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A3_c_315_n N_A_339_368#_c_765_n 0.0113536f $X=4.415 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A3_c_312_n N_A_339_368#_c_785_n 6.60473e-19 $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A3_c_315_n N_A_339_368#_c_785_n 0.0138036f $X=4.415 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A3_c_316_n N_A_339_368#_c_785_n 0.0133547f $X=4.865 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A3_c_317_n N_A_339_368#_c_785_n 6.12174e-19 $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A3_c_311_n N_A_339_368#_c_785_n 0.00124994f $X=5.58 $Y=1.385 $X2=0
+ $Y2=0
cc_302 N_A3_c_316_n N_A_339_368#_c_766_n 0.0108414f $X=4.865 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A3_c_317_n N_A_339_368#_c_766_n 0.0134708f $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A3_c_316_n N_A_339_368#_c_767_n 6.12174e-19 $X=4.865 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A3_c_317_n N_A_339_368#_c_767_n 0.015659f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_306 N_A3_c_312_n N_A_339_368#_c_769_n 0.00171731f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A3_c_315_n N_A_339_368#_c_770_n 0.00175197f $X=4.415 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_A3_c_316_n N_A_339_368#_c_770_n 0.00175197f $X=4.865 $Y=1.765 $X2=0
+ $Y2=0
cc_309 N_A3_c_304_n N_A_788_368#_c_845_n 0.00100811f $X=4.325 $Y=1.65 $X2=0
+ $Y2=0
cc_310 N_A3_c_315_n N_A_788_368#_c_845_n 0.0112044f $X=4.415 $Y=1.765 $X2=0
+ $Y2=0
cc_311 N_A3_c_316_n N_A_788_368#_c_845_n 0.0103758f $X=4.865 $Y=1.765 $X2=0
+ $Y2=0
cc_312 A3 N_A_788_368#_c_845_n 0.0417698f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_313 N_A3_c_311_n N_A_788_368#_c_845_n 0.0206448f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_314 N_A3_c_312_n N_A_788_368#_c_841_n 0.0013314f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_315 N_A3_c_304_n N_A_788_368#_c_841_n 0.015687f $X=4.325 $Y=1.65 $X2=0 $Y2=0
cc_316 N_A3_c_305_n N_A_788_368#_c_841_n 7.51749e-19 $X=3.955 $Y=1.65 $X2=0
+ $Y2=0
cc_317 N_A3_c_317_n N_A_788_368#_c_842_n 0.0117819f $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_318 A3 N_A_788_368#_c_842_n 0.0697636f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_319 N_A3_c_311_n N_A_788_368#_c_842_n 0.0147882f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_320 A3 N_A_788_368#_c_856_n 0.0185129f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_321 N_A3_c_311_n N_A_788_368#_c_856_n 0.00919994f $X=5.58 $Y=1.385 $X2=0
+ $Y2=0
cc_322 N_A3_c_317_n N_A_1191_368#_c_888_n 0.00206065f $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A3_c_317_n N_A_1191_368#_c_890_n 6.23416e-19 $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_A3_c_304_n N_A_27_74#_c_976_n 0.00355178f $X=4.325 $Y=1.65 $X2=0 $Y2=0
cc_325 N_A3_c_305_n N_A_27_74#_c_976_n 0.00449537f $X=3.955 $Y=1.65 $X2=0 $Y2=0
cc_326 A3 N_A_27_74#_c_976_n 0.013152f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_327 N_A3_c_311_n N_A_27_74#_c_976_n 0.00422915f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_328 N_A3_c_306_n N_A_27_74#_c_977_n 0.00722697f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_329 N_A3_c_307_n N_A_27_74#_c_977_n 7.0998e-19 $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_330 N_A3_c_306_n N_A_27_74#_c_978_n 0.00418933f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_331 A3 N_A_27_74#_c_978_n 0.00818182f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_332 N_A3_c_306_n N_A_27_74#_c_1033_n 0.010267f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_333 N_A3_c_307_n N_A_27_74#_c_1033_n 0.0100105f $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_334 A3 N_A_27_74#_c_1033_n 0.0422704f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_335 N_A3_c_311_n N_A_27_74#_c_1033_n 0.00106584f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_336 N_A3_c_307_n N_A_27_74#_c_979_n 2.29136e-19 $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_337 N_A3_c_308_n N_A_27_74#_c_979_n 0.00703259f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_338 N_A3_c_309_n N_A_27_74#_c_979_n 7.13338e-19 $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_339 N_A3_c_308_n N_A_27_74#_c_1040_n 0.00892313f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_340 N_A3_c_309_n N_A_27_74#_c_1040_n 0.0100105f $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_341 A3 N_A_27_74#_c_1040_n 0.0454799f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_342 N_A3_c_311_n N_A_27_74#_c_1040_n 0.00107356f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_343 N_A3_c_309_n N_A_27_74#_c_980_n 2.29136e-19 $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_344 N_A3_c_304_n N_A_27_74#_c_1024_n 0.00272769f $X=4.325 $Y=1.65 $X2=0 $Y2=0
cc_345 N_A3_c_306_n N_A_27_74#_c_1024_n 0.00157416f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_346 N_A3_c_308_n N_A_27_74#_c_1047_n 7.17169e-19 $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_347 A3 N_A_27_74#_c_1047_n 0.0189543f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_348 N_A3_c_311_n N_A_27_74#_c_1047_n 7.01515e-19 $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_349 A3 N_A_27_74#_c_1050_n 0.0134301f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_350 N_A3_c_306_n N_VGND_c_1161_n 0.00434272f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_351 N_A3_c_306_n N_VGND_c_1162_n 0.00482414f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_352 N_A3_c_307_n N_VGND_c_1162_n 0.00771106f $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_353 N_A3_c_308_n N_VGND_c_1162_n 4.39845e-19 $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_354 N_A3_c_307_n N_VGND_c_1163_n 0.00383152f $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_355 N_A3_c_308_n N_VGND_c_1163_n 0.00434272f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_356 N_A3_c_308_n N_VGND_c_1164_n 0.00335277f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_357 N_A3_c_309_n N_VGND_c_1164_n 0.00771106f $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_358 N_A3_c_309_n N_VGND_c_1172_n 0.00383152f $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_359 N_A3_c_306_n N_VGND_c_1177_n 0.00445593f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_360 N_A3_c_307_n N_VGND_c_1177_n 0.00383967f $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_361 N_A3_c_308_n N_VGND_c_1177_n 0.00445496f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_362 N_A3_c_309_n N_VGND_c_1177_n 0.00384065f $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_363 N_A2_c_417_n N_A1_c_509_n 0.0111674f $X=7.675 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_364 N_A2_c_411_n N_A1_c_503_n 0.00901198f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_365 A2 N_A1_c_503_n 0.00453332f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_366 A2 A1 0.0247094f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_367 N_A2_c_413_n A1 2.11798e-19 $X=7.655 $Y=1.492 $X2=0 $Y2=0
cc_368 N_A2_c_413_n N_A1_c_508_n 0.0248291f $X=7.655 $Y=1.492 $X2=0 $Y2=0
cc_369 N_A2_c_417_n N_VPWR_c_585_n 4.40806e-19 $X=7.675 $Y=1.765 $X2=0 $Y2=0
cc_370 N_A2_c_414_n N_VPWR_c_588_n 0.00278257f $X=6.325 $Y=1.765 $X2=0 $Y2=0
cc_371 N_A2_c_415_n N_VPWR_c_588_n 0.00278257f $X=6.775 $Y=1.765 $X2=0 $Y2=0
cc_372 N_A2_c_416_n N_VPWR_c_588_n 0.00278257f $X=7.225 $Y=1.765 $X2=0 $Y2=0
cc_373 N_A2_c_417_n N_VPWR_c_588_n 0.00278257f $X=7.675 $Y=1.765 $X2=0 $Y2=0
cc_374 N_A2_c_414_n N_VPWR_c_581_n 0.00358623f $X=6.325 $Y=1.765 $X2=0 $Y2=0
cc_375 N_A2_c_415_n N_VPWR_c_581_n 0.00353822f $X=6.775 $Y=1.765 $X2=0 $Y2=0
cc_376 N_A2_c_416_n N_VPWR_c_581_n 0.00353822f $X=7.225 $Y=1.765 $X2=0 $Y2=0
cc_377 N_A2_c_417_n N_VPWR_c_581_n 0.00353905f $X=7.675 $Y=1.765 $X2=0 $Y2=0
cc_378 N_A2_c_414_n N_A_339_368#_c_766_n 5.92854e-19 $X=6.325 $Y=1.765 $X2=0
+ $Y2=0
cc_379 N_A2_c_414_n N_A_339_368#_c_767_n 0.00208616f $X=6.325 $Y=1.765 $X2=0
+ $Y2=0
cc_380 N_A2_c_414_n N_A_788_368#_c_842_n 0.0117819f $X=6.325 $Y=1.765 $X2=0
+ $Y2=0
cc_381 A2 N_A_788_368#_c_842_n 0.00508283f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_382 N_A2_c_413_n N_A_788_368#_c_842_n 0.0113335f $X=7.655 $Y=1.492 $X2=0
+ $Y2=0
cc_383 N_A2_c_415_n N_A_788_368#_c_843_n 0.0103384f $X=6.775 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A2_c_416_n N_A_788_368#_c_843_n 0.0103162f $X=7.225 $Y=1.765 $X2=0
+ $Y2=0
cc_385 N_A2_c_417_n N_A_788_368#_c_843_n 6.88765e-19 $X=7.675 $Y=1.765 $X2=0
+ $Y2=0
cc_386 A2 N_A_788_368#_c_843_n 0.0689321f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_387 N_A2_c_413_n N_A_788_368#_c_843_n 0.0139592f $X=7.655 $Y=1.492 $X2=0
+ $Y2=0
cc_388 A2 N_A_788_368#_c_844_n 0.0195526f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_389 N_A2_c_413_n N_A_788_368#_c_844_n 0.00209661f $X=7.655 $Y=1.492 $X2=0
+ $Y2=0
cc_390 N_A2_c_414_n N_A_1191_368#_c_888_n 0.0155173f $X=6.325 $Y=1.765 $X2=0
+ $Y2=0
cc_391 N_A2_c_415_n N_A_1191_368#_c_888_n 6.08256e-19 $X=6.775 $Y=1.765 $X2=0
+ $Y2=0
cc_392 N_A2_c_414_n N_A_1191_368#_c_889_n 0.011279f $X=6.325 $Y=1.765 $X2=0
+ $Y2=0
cc_393 N_A2_c_415_n N_A_1191_368#_c_889_n 0.011279f $X=6.775 $Y=1.765 $X2=0
+ $Y2=0
cc_394 N_A2_c_414_n N_A_1191_368#_c_890_n 0.00264911f $X=6.325 $Y=1.765 $X2=0
+ $Y2=0
cc_395 N_A2_c_414_n N_A_1191_368#_c_906_n 6.08256e-19 $X=6.325 $Y=1.765 $X2=0
+ $Y2=0
cc_396 N_A2_c_415_n N_A_1191_368#_c_906_n 0.0132129f $X=6.775 $Y=1.765 $X2=0
+ $Y2=0
cc_397 N_A2_c_416_n N_A_1191_368#_c_906_n 0.0130919f $X=7.225 $Y=1.765 $X2=0
+ $Y2=0
cc_398 N_A2_c_417_n N_A_1191_368#_c_906_n 5.6787e-19 $X=7.675 $Y=1.765 $X2=0
+ $Y2=0
cc_399 N_A2_c_416_n N_A_1191_368#_c_891_n 0.0107904f $X=7.225 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_A2_c_417_n N_A_1191_368#_c_891_n 0.0123223f $X=7.675 $Y=1.765 $X2=0
+ $Y2=0
cc_401 N_A2_c_416_n N_A_1191_368#_c_912_n 6.57759e-19 $X=7.225 $Y=1.765 $X2=0
+ $Y2=0
cc_402 N_A2_c_417_n N_A_1191_368#_c_912_n 0.0118697f $X=7.675 $Y=1.765 $X2=0
+ $Y2=0
cc_403 A2 N_A_1191_368#_c_892_n 0.00156259f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_404 N_A2_c_417_n N_A_1191_368#_c_893_n 0.00207548f $X=7.675 $Y=1.765 $X2=0
+ $Y2=0
cc_405 A2 N_A_1191_368#_c_893_n 0.0247125f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_406 N_A2_c_413_n N_A_1191_368#_c_893_n 0.00184971f $X=7.655 $Y=1.492 $X2=0
+ $Y2=0
cc_407 N_A2_c_415_n N_A_1191_368#_c_897_n 0.00177174f $X=6.775 $Y=1.765 $X2=0
+ $Y2=0
cc_408 N_A2_c_416_n N_A_1191_368#_c_897_n 0.00201554f $X=7.225 $Y=1.765 $X2=0
+ $Y2=0
cc_409 N_A2_c_408_n N_A_27_74#_c_980_n 0.00703259f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_410 N_A2_c_409_n N_A_27_74#_c_980_n 7.13338e-19 $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_411 N_A2_c_408_n N_A_27_74#_c_1053_n 0.0126582f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_412 N_A2_c_409_n N_A_27_74#_c_1053_n 0.0100105f $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_413 A2 N_A_27_74#_c_1053_n 0.0352336f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_414 N_A2_c_413_n N_A_27_74#_c_1053_n 0.00106692f $X=7.655 $Y=1.492 $X2=0
+ $Y2=0
cc_415 N_A2_c_409_n N_A_27_74#_c_981_n 2.23968e-19 $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_416 N_A2_c_410_n N_A_27_74#_c_981_n 2.23968e-19 $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_417 N_A2_c_410_n N_A_27_74#_c_1059_n 0.00982315f $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_418 N_A2_c_411_n N_A_27_74#_c_1059_n 0.0100509f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_419 A2 N_A_27_74#_c_1059_n 0.046858f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_420 N_A2_c_413_n N_A_27_74#_c_1059_n 8.48385e-19 $X=7.655 $Y=1.492 $X2=0
+ $Y2=0
cc_421 N_A2_c_411_n N_A_27_74#_c_982_n 2.6818e-19 $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_422 N_A2_c_408_n N_A_27_74#_c_1050_n 0.00151008f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_423 A2 N_A_27_74#_c_1065_n 0.0146489f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_424 N_A2_c_413_n N_A_27_74#_c_1065_n 7.03576e-19 $X=7.655 $Y=1.492 $X2=0
+ $Y2=0
cc_425 A2 N_A_27_74#_c_1067_n 0.0205097f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_426 N_A2_c_408_n N_VGND_c_1164_n 4.39845e-19 $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_427 N_A2_c_408_n N_VGND_c_1165_n 0.00335277f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_428 N_A2_c_409_n N_VGND_c_1165_n 0.00759025f $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_429 N_A2_c_410_n N_VGND_c_1165_n 4.20905e-19 $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_430 N_A2_c_409_n N_VGND_c_1166_n 4.20905e-19 $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_431 N_A2_c_410_n N_VGND_c_1166_n 0.00749469f $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_432 N_A2_c_411_n N_VGND_c_1166_n 0.00192221f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_433 N_A2_c_411_n N_VGND_c_1167_n 4.08135e-19 $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_434 N_A2_c_408_n N_VGND_c_1172_n 0.00434272f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_435 N_A2_c_409_n N_VGND_c_1173_n 0.00383152f $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_436 N_A2_c_410_n N_VGND_c_1173_n 0.00383152f $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_437 N_A2_c_411_n N_VGND_c_1174_n 0.00461464f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_438 N_A2_c_408_n N_VGND_c_1177_n 0.00445593f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_439 N_A2_c_409_n N_VGND_c_1177_n 0.00383967f $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_440 N_A2_c_410_n N_VGND_c_1177_n 0.00383967f $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_441 N_A2_c_411_n N_VGND_c_1177_n 0.00463521f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_442 N_A1_c_509_n N_VPWR_c_585_n 0.0143167f $X=8.125 $Y=1.765 $X2=0 $Y2=0
cc_443 N_A1_c_510_n N_VPWR_c_585_n 0.0065594f $X=8.625 $Y=1.765 $X2=0 $Y2=0
cc_444 N_A1_c_511_n N_VPWR_c_586_n 0.0065594f $X=9.075 $Y=1.765 $X2=0 $Y2=0
cc_445 N_A1_c_512_n N_VPWR_c_586_n 0.0175296f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_446 N_A1_c_509_n N_VPWR_c_588_n 0.00413917f $X=8.125 $Y=1.765 $X2=0 $Y2=0
cc_447 N_A1_c_510_n N_VPWR_c_589_n 0.00445347f $X=8.625 $Y=1.765 $X2=0 $Y2=0
cc_448 N_A1_c_511_n N_VPWR_c_589_n 0.00445347f $X=9.075 $Y=1.765 $X2=0 $Y2=0
cc_449 N_A1_c_512_n N_VPWR_c_590_n 0.00413917f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_450 N_A1_c_509_n N_VPWR_c_581_n 0.0081781f $X=8.125 $Y=1.765 $X2=0 $Y2=0
cc_451 N_A1_c_510_n N_VPWR_c_581_n 0.008572f $X=8.625 $Y=1.765 $X2=0 $Y2=0
cc_452 N_A1_c_511_n N_VPWR_c_581_n 0.008572f $X=9.075 $Y=1.765 $X2=0 $Y2=0
cc_453 N_A1_c_512_n N_VPWR_c_581_n 0.00821221f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_454 N_A1_c_509_n N_A_1191_368#_c_891_n 9.96279e-19 $X=8.125 $Y=1.765 $X2=0
+ $Y2=0
cc_455 N_A1_c_509_n N_A_1191_368#_c_892_n 0.0105536f $X=8.125 $Y=1.765 $X2=0
+ $Y2=0
cc_456 N_A1_c_510_n N_A_1191_368#_c_892_n 0.0092358f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_457 A1 N_A_1191_368#_c_892_n 0.0297341f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_458 N_A1_c_508_n N_A_1191_368#_c_892_n 0.0167635f $X=9.575 $Y=1.492 $X2=0
+ $Y2=0
cc_459 N_A1_c_509_n N_A_1191_368#_c_894_n 7.76646e-19 $X=8.125 $Y=1.765 $X2=0
+ $Y2=0
cc_460 N_A1_c_510_n N_A_1191_368#_c_894_n 0.0139897f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_461 N_A1_c_511_n N_A_1191_368#_c_894_n 0.0139897f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_462 N_A1_c_512_n N_A_1191_368#_c_894_n 7.76646e-19 $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_463 N_A1_c_511_n N_A_1191_368#_c_895_n 0.0092358f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_464 N_A1_c_512_n N_A_1191_368#_c_895_n 0.0111377f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_465 A1 N_A_1191_368#_c_895_n 0.0736603f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_466 N_A1_c_508_n N_A_1191_368#_c_895_n 0.0118201f $X=9.575 $Y=1.492 $X2=0
+ $Y2=0
cc_467 N_A1_c_512_n N_A_1191_368#_c_896_n 0.00267251f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_468 N_A1_c_510_n N_A_1191_368#_c_898_n 0.00109449f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_469 N_A1_c_511_n N_A_1191_368#_c_898_n 0.00109449f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_470 A1 N_A_1191_368#_c_898_n 0.0277828f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_471 N_A1_c_508_n N_A_1191_368#_c_898_n 0.00507541f $X=9.575 $Y=1.492 $X2=0
+ $Y2=0
cc_472 N_A1_c_503_n N_A_27_74#_c_982_n 2.68041e-19 $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_473 N_A1_c_503_n N_A_27_74#_c_1069_n 0.0147786f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_474 N_A1_c_504_n N_A_27_74#_c_1069_n 0.00899821f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_475 A1 N_A_27_74#_c_1069_n 0.0301154f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_476 N_A1_c_508_n N_A_27_74#_c_1069_n 0.00116455f $X=9.575 $Y=1.492 $X2=0
+ $Y2=0
cc_477 N_A1_c_503_n N_A_27_74#_c_983_n 4.37256e-19 $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_478 N_A1_c_504_n N_A_27_74#_c_983_n 0.0073734f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_479 N_A1_c_505_n N_A_27_74#_c_983_n 0.00723778f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_480 N_A1_c_506_n N_A_27_74#_c_983_n 7.0998e-19 $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_481 N_A1_c_505_n N_A_27_74#_c_1077_n 0.00892313f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_482 N_A1_c_506_n N_A_27_74#_c_1077_n 0.0100105f $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_483 A1 N_A_27_74#_c_1077_n 0.0454799f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_484 N_A1_c_508_n N_A_27_74#_c_1077_n 0.00107107f $X=9.575 $Y=1.492 $X2=0
+ $Y2=0
cc_485 A1 N_A_27_74#_c_984_n 0.0208616f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_486 N_A1_c_506_n N_A_27_74#_c_985_n 8.26992e-19 $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_487 N_A1_c_504_n N_A_27_74#_c_1083_n 7.17169e-19 $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_488 N_A1_c_505_n N_A_27_74#_c_1083_n 7.17169e-19 $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_489 A1 N_A_27_74#_c_1083_n 0.0232596f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_490 N_A1_c_508_n N_A_27_74#_c_1083_n 7.03992e-19 $X=9.575 $Y=1.492 $X2=0
+ $Y2=0
cc_491 N_A1_c_503_n N_VGND_c_1167_n 0.00685728f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_492 N_A1_c_504_n N_VGND_c_1167_n 0.00352333f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_493 N_A1_c_505_n N_VGND_c_1168_n 0.00344221f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_494 N_A1_c_506_n N_VGND_c_1168_n 0.0105358f $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_495 N_A1_c_503_n N_VGND_c_1174_n 0.00429299f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_496 N_A1_c_504_n N_VGND_c_1175_n 0.00434272f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_497 N_A1_c_505_n N_VGND_c_1175_n 0.00434272f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_498 N_A1_c_506_n N_VGND_c_1176_n 0.00383152f $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_499 N_A1_c_503_n N_VGND_c_1177_n 0.00430064f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_500 N_A1_c_504_n N_VGND_c_1177_n 0.00445625f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_501 N_A1_c_505_n N_VGND_c_1177_n 0.00445496f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_502 N_A1_c_506_n N_VGND_c_1177_n 0.00387625f $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_503 N_VPWR_c_583_n N_Y_c_689_n 0.0416899f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_504 N_VPWR_c_584_n N_Y_c_689_n 0.0353111f $X=1.28 $Y=2.225 $X2=0 $Y2=0
cc_505 N_VPWR_c_587_n N_Y_c_689_n 0.0146357f $X=1.115 $Y=3.33 $X2=0 $Y2=0
cc_506 N_VPWR_c_581_n N_Y_c_689_n 0.0121141f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_507 N_VPWR_M1026_d N_Y_c_690_n 0.0028012f $X=1.13 $Y=1.84 $X2=0 $Y2=0
cc_508 N_VPWR_c_584_n N_Y_c_690_n 0.0219924f $X=1.28 $Y=2.225 $X2=0 $Y2=0
cc_509 N_VPWR_c_583_n N_Y_c_691_n 0.0035248f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_510 N_VPWR_c_584_n N_A_339_368#_c_760_n 0.0565979f $X=1.28 $Y=2.225 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_588_n N_A_339_368#_c_761_n 0.0390078f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_581_n N_A_339_368#_c_761_n 0.0219374f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_584_n N_A_339_368#_c_762_n 0.0121617f $X=1.28 $Y=2.225 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_588_n N_A_339_368#_c_762_n 0.0218645f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_581_n N_A_339_368#_c_762_n 0.0118577f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_588_n N_A_339_368#_c_763_n 0.0390078f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_581_n N_A_339_368#_c_763_n 0.0219374f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_588_n N_A_339_368#_c_765_n 0.0423218f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_581_n N_A_339_368#_c_765_n 0.0239549f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_588_n N_A_339_368#_c_766_n 0.0594839f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_581_n N_A_339_368#_c_766_n 0.0329562f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_588_n N_A_339_368#_c_768_n 0.0200723f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_581_n N_A_339_368#_c_768_n 0.0108858f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_588_n N_A_339_368#_c_769_n 0.0218117f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_581_n N_A_339_368#_c_769_n 0.0117891f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_588_n N_A_339_368#_c_770_n 0.0235512f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_581_n N_A_339_368#_c_770_n 0.0126924f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_588_n N_A_1191_368#_c_889_n 0.0360853f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_581_n N_A_1191_368#_c_889_n 0.0202329f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_588_n N_A_1191_368#_c_890_n 0.0236039f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_581_n N_A_1191_368#_c_890_n 0.012761f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_585_n N_A_1191_368#_c_891_n 0.0117237f $X=8.35 $Y=2.225 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_588_n N_A_1191_368#_c_891_n 0.0558996f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_581_n N_A_1191_368#_c_891_n 0.0310123f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_M1018_s N_A_1191_368#_c_892_n 0.00250873f $X=8.2 $Y=1.84 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_585_n N_A_1191_368#_c_892_n 0.0202249f $X=8.35 $Y=2.225 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_585_n N_A_1191_368#_c_894_n 0.0368936f $X=8.35 $Y=2.225 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_586_n N_A_1191_368#_c_894_n 0.0368936f $X=9.35 $Y=2.225 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_589_n N_A_1191_368#_c_894_n 0.0158233f $X=9.185 $Y=3.33 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_581_n N_A_1191_368#_c_894_n 0.0121241f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_M1020_s N_A_1191_368#_c_895_n 0.00250873f $X=9.15 $Y=1.84 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_586_n N_A_1191_368#_c_895_n 0.0202249f $X=9.35 $Y=2.225 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_586_n N_A_1191_368#_c_896_n 0.0368538f $X=9.35 $Y=2.225 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_590_n N_A_1191_368#_c_896_n 0.0134846f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_581_n N_A_1191_368#_c_896_n 0.0103893f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_588_n N_A_1191_368#_c_897_n 0.0235512f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_581_n N_A_1191_368#_c_897_n 0.0126924f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_Y_c_693_n N_A_339_368#_M1000_s 0.00135003f $X=2.15 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_549 N_Y_c_695_n N_A_339_368#_M1000_s 0.00149404f $X=1.64 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_550 N_Y_c_728_n N_A_339_368#_M1004_s 0.00203444f $X=3.05 $Y=1.935 $X2=0 $Y2=0
cc_551 N_Y_c_693_n N_A_339_368#_c_760_n 0.0103774f $X=2.15 $Y=1.805 $X2=0 $Y2=0
cc_552 N_Y_c_695_n N_A_339_368#_c_760_n 0.011698f $X=1.64 $Y=1.805 $X2=0 $Y2=0
cc_553 N_Y_M1000_d N_A_339_368#_c_761_n 0.00197722f $X=2.14 $Y=1.84 $X2=0 $Y2=0
cc_554 N_Y_c_745_p N_A_339_368#_c_761_n 0.014157f $X=2.29 $Y=2.57 $X2=0 $Y2=0
cc_555 N_Y_c_728_n N_A_339_368#_c_775_n 0.0161421f $X=3.05 $Y=1.935 $X2=0 $Y2=0
cc_556 N_Y_M1029_d N_A_339_368#_c_763_n 0.00197722f $X=3.04 $Y=1.84 $X2=0 $Y2=0
cc_557 N_Y_c_748_p N_A_339_368#_c_763_n 0.014157f $X=3.19 $Y=2.57 $X2=0 $Y2=0
cc_558 N_Y_c_694_n N_A_339_368#_c_764_n 0.00342816f $X=3.19 $Y=2.15 $X2=0 $Y2=0
cc_559 N_Y_c_694_n N_A_788_368#_c_841_n 0.002673f $X=3.19 $Y=2.15 $X2=0 $Y2=0
cc_560 N_Y_c_698_n N_A_27_74#_M1022_d 0.00433624f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_561 N_Y_M1017_s N_A_27_74#_c_971_n 0.00176461f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_562 N_Y_c_698_n N_A_27_74#_c_971_n 0.0035136f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_563 N_Y_c_715_n N_A_27_74#_c_971_n 0.0121701f $X=0.71 $Y=0.8 $X2=0 $Y2=0
cc_564 N_Y_M1030_s N_A_27_74#_c_973_n 0.00250873f $X=1.43 $Y=0.37 $X2=0 $Y2=0
cc_565 N_Y_c_698_n N_A_27_74#_c_973_n 0.00352531f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_566 N_Y_c_708_n N_A_27_74#_c_973_n 0.019744f $X=1.64 $Y=1.01 $X2=0 $Y2=0
cc_567 N_Y_c_698_n N_A_27_74#_c_986_n 0.0160355f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_568 N_Y_c_698_n N_VGND_c_1177_n 0.00143802f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_569 N_A_339_368#_c_765_n N_A_788_368#_M1001_s 0.00315979f $X=4.475 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_570 N_A_339_368#_c_766_n N_A_788_368#_M1007_s 0.00197722f $X=5.375 $Y=2.99
+ $X2=0 $Y2=0
cc_571 N_A_339_368#_c_765_n N_A_788_368#_c_871_n 0.0217683f $X=4.475 $Y=2.99
+ $X2=0 $Y2=0
cc_572 N_A_339_368#_M1006_d N_A_788_368#_c_845_n 0.00197722f $X=4.49 $Y=1.84
+ $X2=0 $Y2=0
cc_573 N_A_339_368#_c_785_n N_A_788_368#_c_845_n 0.0171813f $X=4.64 $Y=2.145
+ $X2=0 $Y2=0
cc_574 N_A_339_368#_c_764_n N_A_788_368#_c_841_n 0.00517051f $X=3.64 $Y=1.965
+ $X2=0 $Y2=0
cc_575 N_A_339_368#_c_766_n N_A_788_368#_c_875_n 0.014157f $X=5.375 $Y=2.99
+ $X2=0 $Y2=0
cc_576 N_A_339_368#_M1014_d N_A_788_368#_c_842_n 0.0028012f $X=5.39 $Y=1.84
+ $X2=0 $Y2=0
cc_577 N_A_339_368#_c_767_n N_A_788_368#_c_842_n 0.0219924f $X=5.54 $Y=2.145
+ $X2=0 $Y2=0
cc_578 N_A_339_368#_c_767_n N_A_1191_368#_c_888_n 0.0559238f $X=5.54 $Y=2.145
+ $X2=0 $Y2=0
cc_579 N_A_339_368#_c_766_n N_A_1191_368#_c_890_n 0.0128665f $X=5.375 $Y=2.99
+ $X2=0 $Y2=0
cc_580 N_A_339_368#_c_767_n N_A_1191_368#_c_890_n 0.00103928f $X=5.54 $Y=2.145
+ $X2=0 $Y2=0
cc_581 N_A_339_368#_c_764_n N_A_27_74#_c_976_n 0.01605f $X=3.64 $Y=1.965 $X2=0
+ $Y2=0
cc_582 N_A_788_368#_c_842_n N_A_1191_368#_M1009_s 0.0028012f $X=6.435 $Y=1.805
+ $X2=-0.19 $Y2=1.66
cc_583 N_A_788_368#_c_843_n N_A_1191_368#_M1010_s 0.00197722f $X=7.335 $Y=1.805
+ $X2=0 $Y2=0
cc_584 N_A_788_368#_c_842_n N_A_1191_368#_c_888_n 0.0219924f $X=6.435 $Y=1.805
+ $X2=0 $Y2=0
cc_585 N_A_788_368#_M1009_d N_A_1191_368#_c_889_n 0.00198238f $X=6.4 $Y=1.84
+ $X2=0 $Y2=0
cc_586 N_A_788_368#_c_882_p N_A_1191_368#_c_889_n 0.0142892f $X=6.55 $Y=1.965
+ $X2=0 $Y2=0
cc_587 N_A_788_368#_c_843_n N_A_1191_368#_c_906_n 0.0171813f $X=7.335 $Y=1.805
+ $X2=0 $Y2=0
cc_588 N_A_788_368#_M1013_d N_A_1191_368#_c_891_n 0.00197722f $X=7.3 $Y=1.84
+ $X2=0 $Y2=0
cc_589 N_A_788_368#_c_885_p N_A_1191_368#_c_891_n 0.014157f $X=7.45 $Y=2.045
+ $X2=0 $Y2=0
cc_590 N_A_788_368#_c_843_n N_A_1191_368#_c_893_n 0.012724f $X=7.335 $Y=1.805
+ $X2=0 $Y2=0
cc_591 N_A_788_368#_c_841_n N_A_27_74#_c_976_n 0.0139914f $X=4.305 $Y=1.805
+ $X2=0 $Y2=0
cc_592 N_A_27_74#_c_1002_n N_VGND_M1002_d 0.0117286f $X=3.16 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_593 N_A_27_74#_c_1033_n N_VGND_M1003_d 0.00462121f $X=5.03 $Y=0.925 $X2=0
+ $Y2=0
cc_594 N_A_27_74#_c_1040_n N_VGND_M1036_d 0.00462121f $X=5.96 $Y=0.925 $X2=0
+ $Y2=0
cc_595 N_A_27_74#_c_1053_n N_VGND_M1005_s 0.00462121f $X=6.89 $Y=0.925 $X2=0
+ $Y2=0
cc_596 N_A_27_74#_c_1059_n N_VGND_M1025_s 0.00395707f $X=7.785 $Y=0.925 $X2=0
+ $Y2=0
cc_597 N_A_27_74#_c_1069_n N_VGND_M1008_s 0.00530982f $X=8.705 $Y=0.925 $X2=0
+ $Y2=0
cc_598 N_A_27_74#_c_1077_n N_VGND_M1033_s 0.00462121f $X=9.715 $Y=0.925 $X2=0
+ $Y2=0
cc_599 N_A_27_74#_c_974_n N_VGND_c_1160_n 0.0191473f $X=3.325 $Y=0.515 $X2=0
+ $Y2=0
cc_600 N_A_27_74#_c_975_n N_VGND_c_1160_n 0.00474779f $X=3.415 $Y=1.3 $X2=0
+ $Y2=0
cc_601 N_A_27_74#_c_976_n N_VGND_c_1160_n 0.013555f $X=4.02 $Y=1.385 $X2=0 $Y2=0
cc_602 N_A_27_74#_c_977_n N_VGND_c_1160_n 0.018213f $X=4.185 $Y=0.515 $X2=0
+ $Y2=0
cc_603 N_A_27_74#_c_978_n N_VGND_c_1160_n 0.00453882f $X=4.105 $Y=1.3 $X2=0
+ $Y2=0
cc_604 N_A_27_74#_c_977_n N_VGND_c_1161_n 0.014477f $X=4.185 $Y=0.515 $X2=0
+ $Y2=0
cc_605 N_A_27_74#_c_977_n N_VGND_c_1162_n 0.0127977f $X=4.185 $Y=0.515 $X2=0
+ $Y2=0
cc_606 N_A_27_74#_c_1033_n N_VGND_c_1162_n 0.0205261f $X=5.03 $Y=0.925 $X2=0
+ $Y2=0
cc_607 N_A_27_74#_c_979_n N_VGND_c_1162_n 0.0121972f $X=5.115 $Y=0.515 $X2=0
+ $Y2=0
cc_608 N_A_27_74#_c_979_n N_VGND_c_1163_n 0.0109704f $X=5.115 $Y=0.515 $X2=0
+ $Y2=0
cc_609 N_A_27_74#_c_979_n N_VGND_c_1164_n 0.0122975f $X=5.115 $Y=0.515 $X2=0
+ $Y2=0
cc_610 N_A_27_74#_c_1040_n N_VGND_c_1164_n 0.0205261f $X=5.96 $Y=0.925 $X2=0
+ $Y2=0
cc_611 N_A_27_74#_c_980_n N_VGND_c_1164_n 0.0121972f $X=6.045 $Y=0.515 $X2=0
+ $Y2=0
cc_612 N_A_27_74#_c_980_n N_VGND_c_1165_n 0.0122975f $X=6.045 $Y=0.515 $X2=0
+ $Y2=0
cc_613 N_A_27_74#_c_1053_n N_VGND_c_1165_n 0.0205261f $X=6.89 $Y=0.925 $X2=0
+ $Y2=0
cc_614 N_A_27_74#_c_981_n N_VGND_c_1165_n 0.0121558f $X=6.975 $Y=0.515 $X2=0
+ $Y2=0
cc_615 N_A_27_74#_c_981_n N_VGND_c_1166_n 0.0121558f $X=6.975 $Y=0.515 $X2=0
+ $Y2=0
cc_616 N_A_27_74#_c_1059_n N_VGND_c_1166_n 0.0177409f $X=7.785 $Y=0.925 $X2=0
+ $Y2=0
cc_617 N_A_27_74#_c_982_n N_VGND_c_1166_n 0.00131301f $X=7.87 $Y=0.515 $X2=0
+ $Y2=0
cc_618 N_A_27_74#_c_982_n N_VGND_c_1167_n 0.0127651f $X=7.87 $Y=0.515 $X2=0
+ $Y2=0
cc_619 N_A_27_74#_c_1069_n N_VGND_c_1167_n 0.020602f $X=8.705 $Y=0.925 $X2=0
+ $Y2=0
cc_620 N_A_27_74#_c_983_n N_VGND_c_1167_n 0.0127977f $X=8.87 $Y=0.515 $X2=0
+ $Y2=0
cc_621 N_A_27_74#_c_983_n N_VGND_c_1168_n 0.0127977f $X=8.87 $Y=0.515 $X2=0
+ $Y2=0
cc_622 N_A_27_74#_c_1077_n N_VGND_c_1168_n 0.0205261f $X=9.715 $Y=0.925 $X2=0
+ $Y2=0
cc_623 N_A_27_74#_c_985_n N_VGND_c_1168_n 0.0121972f $X=9.8 $Y=0.515 $X2=0 $Y2=0
cc_624 N_A_27_74#_c_974_n N_VGND_c_1169_n 0.0149638f $X=3.325 $Y=0.515 $X2=0
+ $Y2=0
cc_625 N_A_27_74#_c_971_n N_VGND_c_1171_n 0.0333877f $X=0.975 $Y=0.34 $X2=0
+ $Y2=0
cc_626 N_A_27_74#_c_972_n N_VGND_c_1171_n 0.0235688f $X=0.445 $Y=0.34 $X2=0
+ $Y2=0
cc_627 N_A_27_74#_c_973_n N_VGND_c_1171_n 0.0781546f $X=1.975 $Y=0.34 $X2=0
+ $Y2=0
cc_628 N_A_27_74#_c_1002_n N_VGND_c_1171_n 0.0278307f $X=3.16 $Y=0.925 $X2=0
+ $Y2=0
cc_629 N_A_27_74#_c_974_n N_VGND_c_1171_n 0.0112517f $X=3.325 $Y=0.515 $X2=0
+ $Y2=0
cc_630 N_A_27_74#_c_986_n N_VGND_c_1171_n 0.0225055f $X=1.14 $Y=0.34 $X2=0 $Y2=0
cc_631 N_A_27_74#_c_980_n N_VGND_c_1172_n 0.0109704f $X=6.045 $Y=0.515 $X2=0
+ $Y2=0
cc_632 N_A_27_74#_c_981_n N_VGND_c_1173_n 0.00747999f $X=6.975 $Y=0.515 $X2=0
+ $Y2=0
cc_633 N_A_27_74#_c_982_n N_VGND_c_1174_n 0.0110419f $X=7.87 $Y=0.515 $X2=0
+ $Y2=0
cc_634 N_A_27_74#_c_983_n N_VGND_c_1175_n 0.0144609f $X=8.87 $Y=0.515 $X2=0
+ $Y2=0
cc_635 N_A_27_74#_c_985_n N_VGND_c_1176_n 0.0110419f $X=9.8 $Y=0.515 $X2=0 $Y2=0
cc_636 N_A_27_74#_c_971_n N_VGND_c_1177_n 0.0187857f $X=0.975 $Y=0.34 $X2=0
+ $Y2=0
cc_637 N_A_27_74#_c_972_n N_VGND_c_1177_n 0.0127152f $X=0.445 $Y=0.34 $X2=0
+ $Y2=0
cc_638 N_A_27_74#_c_973_n N_VGND_c_1177_n 0.0366503f $X=1.975 $Y=0.34 $X2=0
+ $Y2=0
cc_639 N_A_27_74#_c_1002_n N_VGND_c_1177_n 0.0117436f $X=3.16 $Y=0.925 $X2=0
+ $Y2=0
cc_640 N_A_27_74#_c_974_n N_VGND_c_1177_n 0.0123131f $X=3.325 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_A_27_74#_c_977_n N_VGND_c_1177_n 0.0118767f $X=4.185 $Y=0.515 $X2=0
+ $Y2=0
cc_642 N_A_27_74#_c_1033_n N_VGND_c_1177_n 0.0113542f $X=5.03 $Y=0.925 $X2=0
+ $Y2=0
cc_643 N_A_27_74#_c_979_n N_VGND_c_1177_n 0.00903439f $X=5.115 $Y=0.515 $X2=0
+ $Y2=0
cc_644 N_A_27_74#_c_1040_n N_VGND_c_1177_n 0.0113542f $X=5.96 $Y=0.925 $X2=0
+ $Y2=0
cc_645 N_A_27_74#_c_980_n N_VGND_c_1177_n 0.00903439f $X=6.045 $Y=0.515 $X2=0
+ $Y2=0
cc_646 N_A_27_74#_c_1053_n N_VGND_c_1177_n 0.0113542f $X=6.89 $Y=0.925 $X2=0
+ $Y2=0
cc_647 N_A_27_74#_c_981_n N_VGND_c_1177_n 0.00619848f $X=6.975 $Y=0.515 $X2=0
+ $Y2=0
cc_648 N_A_27_74#_c_1059_n N_VGND_c_1177_n 0.0126991f $X=7.785 $Y=0.925 $X2=0
+ $Y2=0
cc_649 N_A_27_74#_c_982_n N_VGND_c_1177_n 0.00915013f $X=7.87 $Y=0.515 $X2=0
+ $Y2=0
cc_650 N_A_27_74#_c_1069_n N_VGND_c_1177_n 0.0109057f $X=8.705 $Y=0.925 $X2=0
+ $Y2=0
cc_651 N_A_27_74#_c_983_n N_VGND_c_1177_n 0.0118703f $X=8.87 $Y=0.515 $X2=0
+ $Y2=0
cc_652 N_A_27_74#_c_1077_n N_VGND_c_1177_n 0.0113542f $X=9.715 $Y=0.925 $X2=0
+ $Y2=0
cc_653 N_A_27_74#_c_985_n N_VGND_c_1177_n 0.00915013f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_654 N_A_27_74#_c_986_n N_VGND_c_1177_n 0.0123739f $X=1.14 $Y=0.34 $X2=0 $Y2=0
