* File: sky130_fd_sc_hs__buf_1.pxi.spice
* Created: Thu Aug 27 20:34:19 2020
* 
x_PM_SKY130_FD_SC_HS__BUF_1%A N_A_M1002_g N_A_c_37_n N_A_M1001_g N_A_c_38_n A A
+ PM_SKY130_FD_SC_HS__BUF_1%A
x_PM_SKY130_FD_SC_HS__BUF_1%A_27_164# N_A_27_164#_M1002_s N_A_27_164#_M1001_s
+ N_A_27_164#_c_70_n N_A_27_164#_M1000_g N_A_27_164#_M1003_g N_A_27_164#_c_77_n
+ N_A_27_164#_c_72_n N_A_27_164#_c_78_n N_A_27_164#_c_79_n N_A_27_164#_c_73_n
+ N_A_27_164#_c_74_n N_A_27_164#_c_75_n PM_SKY130_FD_SC_HS__BUF_1%A_27_164#
x_PM_SKY130_FD_SC_HS__BUF_1%VPWR N_VPWR_M1001_d N_VPWR_c_129_n VPWR
+ N_VPWR_c_130_n N_VPWR_c_131_n N_VPWR_c_128_n N_VPWR_c_133_n
+ PM_SKY130_FD_SC_HS__BUF_1%VPWR
x_PM_SKY130_FD_SC_HS__BUF_1%X N_X_M1003_d N_X_M1000_d N_X_c_149_n N_X_c_150_n X
+ X X X N_X_c_151_n PM_SKY130_FD_SC_HS__BUF_1%X
x_PM_SKY130_FD_SC_HS__BUF_1%VGND N_VGND_M1002_d N_VGND_c_174_n VGND
+ N_VGND_c_175_n N_VGND_c_176_n N_VGND_c_177_n N_VGND_c_178_n
+ PM_SKY130_FD_SC_HS__BUF_1%VGND
cc_1 VNB N_A_M1002_g 0.0400717f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.835
cc_2 VNB N_A_c_37_n 0.00733759f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.045
cc_3 VNB N_A_c_38_n 0.0305395f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.615
cc_4 VNB A 0.00958066f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_5 VNB N_A_27_164#_c_70_n 0.0356016f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.54
cc_6 VNB N_A_27_164#_M1003_g 0.0286459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_164#_c_72_n 0.00640208f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_8 VNB N_A_27_164#_c_73_n 0.00728026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_164#_c_74_n 4.08398e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_164#_c_75_n 0.0351504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_VPWR_c_128_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_12 VNB N_X_c_149_n 0.0265168f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.615
cc_13 VNB N_X_c_150_n 0.0135379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_X_c_151_n 0.0246612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_174_n 0.0169218f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.54
cc_16 VNB N_VGND_c_175_n 0.0331697f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_VGND_c_176_n 0.0189562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_177_n 0.146496f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_19 VNB N_VGND_c_178_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_20 VPB N_A_c_37_n 0.0480338f $X=-0.19 $Y=1.66 $X2=0.86 $Y2=2.045
cc_21 VPB N_A_c_38_n 0.0290939f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.615
cc_22 VPB A 0.00913245f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_23 VPB N_A_27_164#_c_70_n 0.0294843f $X=-0.19 $Y=1.66 $X2=0.86 $Y2=2.54
cc_24 VPB N_A_27_164#_c_77_n 0.035396f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.615
cc_25 VPB N_A_27_164#_c_78_n 0.00396888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_26 VPB N_A_27_164#_c_79_n 0.00948019f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_27 VPB N_A_27_164#_c_74_n 0.00295045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_129_n 0.00970163f $X=-0.19 $Y=1.66 $X2=0.86 $Y2=2.54
cc_29 VPB N_VPWR_c_130_n 0.0304483f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_30 VPB N_VPWR_c_131_n 0.0190763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_128_n 0.0671143f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_32 VPB N_VPWR_c_133_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_33 VPB X 0.0138461f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.615
cc_34 VPB X 0.041687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_X_c_151_n 0.00756337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 N_A_M1002_g N_A_27_164#_c_70_n 0.0175909f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_37 N_A_c_37_n N_A_27_164#_c_70_n 0.0323642f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_38 A N_A_27_164#_c_70_n 2.10849e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_39 N_A_M1002_g N_A_27_164#_M1003_g 0.0174961f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_40 N_A_c_37_n N_A_27_164#_c_77_n 0.0137291f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_41 N_A_M1002_g N_A_27_164#_c_72_n 0.0116849f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_42 N_A_c_37_n N_A_27_164#_c_72_n 5.09057e-19 $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_43 N_A_c_37_n N_A_27_164#_c_78_n 0.0130175f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_44 A N_A_27_164#_c_78_n 0.00782149f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_45 N_A_c_37_n N_A_27_164#_c_79_n 0.00458273f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_46 N_A_c_38_n N_A_27_164#_c_79_n 0.00696845f $X=0.77 $Y=1.615 $X2=0 $Y2=0
cc_47 A N_A_27_164#_c_79_n 0.027657f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_48 N_A_M1002_g N_A_27_164#_c_73_n 0.00504032f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_49 A N_A_27_164#_c_73_n 0.0124978f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_50 N_A_c_37_n N_A_27_164#_c_74_n 0.00489705f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_51 A N_A_27_164#_c_74_n 0.00976617f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_52 N_A_M1002_g N_A_27_164#_c_75_n 0.0105457f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_53 N_A_c_38_n N_A_27_164#_c_75_n 0.0121759f $X=0.77 $Y=1.615 $X2=0 $Y2=0
cc_54 A N_A_27_164#_c_75_n 0.0631563f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_55 N_A_c_37_n N_VPWR_c_129_n 0.00737447f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_56 N_A_c_37_n N_VPWR_c_130_n 0.00445602f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_57 N_A_c_37_n N_VPWR_c_128_n 0.00862626f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_58 N_A_M1002_g N_X_c_149_n 8.70516e-19 $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_59 N_A_c_37_n X 7.14264e-19 $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_VGND_c_174_n 0.0060489f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_VGND_c_175_n 0.00451272f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_62 N_A_M1002_g N_VGND_c_177_n 0.00487769f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_63 N_A_27_164#_c_78_n N_VPWR_M1001_d 0.00482878f $X=1.13 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_64 N_A_27_164#_c_74_n N_VPWR_M1001_d 0.00216738f $X=1.215 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_65 N_A_27_164#_c_70_n N_VPWR_c_129_n 0.00776766f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_66 N_A_27_164#_c_77_n N_VPWR_c_129_n 0.0266809f $X=0.635 $Y=2.265 $X2=0 $Y2=0
cc_67 N_A_27_164#_c_78_n N_VPWR_c_129_n 0.0253877f $X=1.13 $Y=2.035 $X2=0 $Y2=0
cc_68 N_A_27_164#_c_77_n N_VPWR_c_130_n 0.0145938f $X=0.635 $Y=2.265 $X2=0 $Y2=0
cc_69 N_A_27_164#_c_70_n N_VPWR_c_131_n 0.00445602f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A_27_164#_c_70_n N_VPWR_c_128_n 0.00861336f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A_27_164#_c_77_n N_VPWR_c_128_n 0.0120466f $X=0.635 $Y=2.265 $X2=0 $Y2=0
cc_72 N_A_27_164#_M1003_g N_X_c_149_n 0.00823464f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A_27_164#_M1003_g N_X_c_150_n 0.00453721f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_27_164#_c_73_n N_X_c_150_n 0.00278159f $X=1.215 $Y=1.63 $X2=0 $Y2=0
cc_75 N_A_27_164#_c_70_n X 0.00303505f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_27_164#_c_73_n X 0.001416f $X=1.215 $Y=1.63 $X2=0 $Y2=0
cc_77 N_A_27_164#_c_74_n X 0.00565815f $X=1.215 $Y=1.95 $X2=0 $Y2=0
cc_78 N_A_27_164#_c_70_n X 0.0126613f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_27_164#_c_77_n X 0.00406709f $X=0.635 $Y=2.265 $X2=0 $Y2=0
cc_80 N_A_27_164#_M1003_g N_X_c_151_n 0.0130801f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_27_164#_c_73_n N_X_c_151_n 0.0309827f $X=1.215 $Y=1.63 $X2=0 $Y2=0
cc_82 N_A_27_164#_c_74_n N_X_c_151_n 0.00622924f $X=1.215 $Y=1.95 $X2=0 $Y2=0
cc_83 N_A_27_164#_c_73_n N_VGND_M1002_d 0.00188126f $X=1.215 $Y=1.63 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_27_164#_c_70_n N_VGND_c_174_n 6.97737e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_27_164#_M1003_g N_VGND_c_174_n 0.00941074f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_86 N_A_27_164#_c_72_n N_VGND_c_174_n 0.0126515f $X=1.13 $Y=1.195 $X2=0 $Y2=0
cc_87 N_A_27_164#_c_73_n N_VGND_c_174_n 0.0150119f $X=1.215 $Y=1.63 $X2=0 $Y2=0
cc_88 N_A_27_164#_M1003_g N_VGND_c_176_n 0.00434272f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_89 N_A_27_164#_M1003_g N_VGND_c_177_n 0.00828717f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_90 N_A_27_164#_c_75_n N_VGND_c_177_n 0.0266705f $X=0.795 $Y=1.04 $X2=0 $Y2=0
cc_91 N_VPWR_c_129_n X 0.027028f $X=1.135 $Y=2.455 $X2=0 $Y2=0
cc_92 N_VPWR_c_131_n X 0.0159324f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_93 N_VPWR_c_128_n X 0.0131546f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_94 N_X_c_149_n N_VGND_c_174_n 0.0231775f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_95 N_X_c_149_n N_VGND_c_176_n 0.0156794f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_96 N_X_c_149_n N_VGND_c_177_n 0.0129217f $X=1.64 $Y=0.515 $X2=0 $Y2=0
