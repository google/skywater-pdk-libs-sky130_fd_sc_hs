* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_27_74# a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_258_392# a_309_338# a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_83_260# a_315_54# a_484_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X3 a_267_80# a_315_54# a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VGND CLK a_984_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_987_393# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 a_477_124# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_315_54# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X8 VGND GATE a_267_80# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_484_508# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X10 VPWR GATE a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X11 VGND a_315_54# a_309_338# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR CLK a_987_393# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X13 a_984_125# a_27_74# a_987_393# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 VPWR a_315_54# a_309_338# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 a_83_260# a_309_338# a_477_124# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 VPWR a_987_393# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X17 a_27_74# a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VGND a_987_393# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_315_54# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
