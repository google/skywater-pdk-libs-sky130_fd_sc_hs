* File: sky130_fd_sc_hs__a2bb2oi_4.pex.spice
* Created: Tue Sep  1 19:52:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%A2_N 1 3 4 6 7 8 9 11 12 13 14 20
c51 4 0 1.88367e-19 $X=0.945 $Y=1.885
r52 27 28 40.0185 $w=5.42e-07 $l=4.5e-07 $layer=POLY_cond $X=0.495 $Y=1.535
+ $X2=0.945 $Y2=1.535
r53 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=1.605 $X2=0.29 $Y2=1.605
r54 18 27 13.7841 $w=5.42e-07 $l=1.55e-07 $layer=POLY_cond $X=0.34 $Y=1.535
+ $X2=0.495 $Y2=1.535
r55 18 24 4.44649 $w=5.42e-07 $l=5e-08 $layer=POLY_cond $X=0.34 $Y=1.535
+ $X2=0.29 $Y2=1.535
r56 18 20 91.1834 $w=4.3e-07 $l=7.05e-07 $layer=POLY_cond $X=0.34 $Y=1.29
+ $X2=0.34 $Y2=0.585
r57 14 25 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.605
r58 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.925
+ $X2=0.29 $Y2=1.295
r59 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.555
+ $X2=0.29 $Y2=0.925
r60 12 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=0.585 $X2=0.29 $Y2=0.585
r61 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.32 $Y=1.185
+ $X2=1.32 $Y2=0.74
r62 8 28 36.3588 $w=5.42e-07 $l=3.1682e-07 $layer=POLY_cond $X=1.035 $Y=1.26
+ $X2=0.945 $Y2=1.535
r63 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.245 $Y=1.26
+ $X2=1.32 $Y2=1.185
r64 7 8 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.245 $Y=1.26
+ $X2=1.035 $Y2=1.26
r65 4 28 33.4577 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.945 $Y=1.885
+ $X2=0.945 $Y2=1.535
r66 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.945 $Y=1.885
+ $X2=0.945 $Y2=2.46
r67 1 27 33.4577 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.495 $Y=1.885
+ $X2=0.495 $Y2=1.535
r68 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.885
+ $X2=0.495 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%A1_N 1 3 6 8 10 11 12 18
c48 18 0 6.19774e-20 $X=1.77 $Y=1.635
c49 6 0 3.63668e-19 $X=1.75 $Y=0.74
r50 18 20 12.3801 $w=2.92e-07 $l=7.5e-08 $layer=POLY_cond $X=1.77 $Y=1.677
+ $X2=1.845 $Y2=1.677
r51 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.635 $X2=1.77 $Y2=1.635
r52 16 18 3.30137 $w=2.92e-07 $l=2e-08 $layer=POLY_cond $X=1.75 $Y=1.677
+ $X2=1.77 $Y2=1.677
r53 15 16 58.5993 $w=2.92e-07 $l=3.55e-07 $layer=POLY_cond $X=1.395 $Y=1.677
+ $X2=1.75 $Y2=1.677
r54 12 19 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.16 $Y=1.635
+ $X2=1.77 $Y2=1.635
r55 11 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.635 $X2=1.77
+ $Y2=1.635
r56 8 20 18.3338 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.845 $Y=1.885
+ $X2=1.845 $Y2=1.677
r57 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.845 $Y=1.885
+ $X2=1.845 $Y2=2.46
r58 4 16 18.3338 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.75 $Y=1.47
+ $X2=1.75 $Y2=1.677
r59 4 6 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.75 $Y=1.47 $X2=1.75
+ $Y2=0.74
r60 1 15 18.3338 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.395 $Y=1.885
+ $X2=1.395 $Y2=1.677
r61 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.395 $Y=1.885
+ $X2=1.395 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%A_114_392# 1 2 7 9 10 11 12 14 15 17 18 20
+ 21 23 24 26 27 28 29 31 32 34 36 37 39 43 45 46 49 53 55 58 62
c150 53 0 6.19774e-20 $X=2.995 $Y=1.34
c151 37 0 1.59797e-19 $X=3.945 $Y=1.475
c152 29 0 9.74273e-21 $X=3.945 $Y=1.765
c153 24 0 1.39795e-19 $X=3.51 $Y=1.22
c154 18 0 1.39795e-19 $X=3.08 $Y=1.22
c155 12 0 1.44963e-19 $X=2.65 $Y=1.22
r156 68 69 1.78079 $w=4.06e-07 $l=1.5e-08 $layer=POLY_cond $X=3.495 $Y=1.492
+ $X2=3.51 $Y2=1.492
r157 65 66 4.15517 $w=4.06e-07 $l=3.5e-08 $layer=POLY_cond $X=3.045 $Y=1.492
+ $X2=3.08 $Y2=1.492
r158 61 65 36.2094 $w=4.06e-07 $l=3.05e-07 $layer=POLY_cond $X=2.74 $Y=1.492
+ $X2=3.045 $Y2=1.492
r159 61 63 10.6847 $w=4.06e-07 $l=9e-08 $layer=POLY_cond $X=2.74 $Y=1.492
+ $X2=2.65 $Y2=1.492
r160 60 62 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=1.34
+ $X2=2.575 $Y2=1.34
r161 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.385 $X2=2.74 $Y2=1.385
r162 56 68 8.90394 $w=4.06e-07 $l=7.5e-08 $layer=POLY_cond $X=3.42 $Y=1.492
+ $X2=3.495 $Y2=1.492
r163 56 66 40.3645 $w=4.06e-07 $l=3.4e-07 $layer=POLY_cond $X=3.42 $Y=1.492
+ $X2=3.08 $Y2=1.492
r164 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.385 $X2=3.42 $Y2=1.385
r165 53 60 6.99698 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=2.995 $Y=1.34
+ $X2=2.74 $Y2=1.34
r166 53 55 11.6616 $w=4.18e-07 $l=4.25e-07 $layer=LI1_cond $X=2.995 $Y=1.34
+ $X2=3.42 $Y2=1.34
r167 52 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=1.215
+ $X2=1.535 $Y2=1.215
r168 52 62 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.62 $Y=1.215
+ $X2=2.575 $Y2=1.215
r169 47 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=1.13
+ $X2=1.535 $Y2=1.215
r170 47 49 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.535 $Y=1.13
+ $X2=1.535 $Y2=0.515
r171 45 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=1.215
+ $X2=1.535 $Y2=1.215
r172 45 46 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.45 $Y=1.215
+ $X2=0.885 $Y2=1.215
r173 41 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.76 $Y=1.3
+ $X2=0.885 $Y2=1.215
r174 41 43 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=0.76 $Y=1.3
+ $X2=0.76 $Y2=2.105
r175 34 39 114.876 $w=1.8e-07 $l=2.9e-07 $layer=POLY_cond $X=4.395 $Y=1.765
+ $X2=4.395 $Y2=1.475
r176 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.395 $Y=1.765
+ $X2=4.395 $Y2=2.4
r177 33 37 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.035 $Y=1.475
+ $X2=3.945 $Y2=1.475
r178 32 39 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.305 $Y=1.475
+ $X2=4.395 $Y2=1.475
r179 32 33 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.305 $Y=1.475
+ $X2=4.035 $Y2=1.475
r180 29 37 114.876 $w=1.8e-07 $l=2.9e-07 $layer=POLY_cond $X=3.945 $Y=1.765
+ $X2=3.945 $Y2=1.475
r181 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.945 $Y=1.765
+ $X2=3.945 $Y2=2.4
r182 28 69 29.0202 $w=4.06e-07 $l=8.30662e-08 $layer=POLY_cond $X=3.585 $Y=1.475
+ $X2=3.51 $Y2=1.492
r183 27 37 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=1.475
+ $X2=3.945 $Y2=1.475
r184 27 28 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.855 $Y=1.475
+ $X2=3.585 $Y2=1.475
r185 24 69 26.2263 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.51 $Y=1.22
+ $X2=3.51 $Y2=1.492
r186 24 26 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.51 $Y=1.22
+ $X2=3.51 $Y2=0.74
r187 21 68 26.2263 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.495 $Y=1.765
+ $X2=3.495 $Y2=1.492
r188 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.495 $Y=1.765
+ $X2=3.495 $Y2=2.4
r189 18 66 26.2263 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.08 $Y=1.22
+ $X2=3.08 $Y2=1.492
r190 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.08 $Y=1.22
+ $X2=3.08 $Y2=0.74
r191 15 65 26.2263 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.045 $Y=1.765
+ $X2=3.045 $Y2=1.492
r192 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.045 $Y=1.765
+ $X2=3.045 $Y2=2.4
r193 12 63 26.2263 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.65 $Y=1.22
+ $X2=2.65 $Y2=1.492
r194 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.65 $Y=1.22
+ $X2=2.65 $Y2=0.74
r195 10 63 29.0202 $w=4.06e-07 $l=2.31482e-07 $layer=POLY_cond $X=2.575 $Y=1.295
+ $X2=2.65 $Y2=1.492
r196 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.575 $Y=1.295
+ $X2=2.295 $Y2=1.295
r197 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.22 $Y=1.22
+ $X2=2.295 $Y2=1.295
r198 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.22 $Y=1.22 $X2=2.22
+ $Y2=0.74
r199 2 43 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.96 $X2=0.72 $Y2=2.105
r200 1 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.395
+ $Y=0.37 $X2=1.535 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 32 49
c85 32 0 1.6954e-19 $X=6 $Y=1.665
r86 49 50 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=6.195 $Y=1.557
+ $X2=6.2 $Y2=1.557
r87 47 49 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=5.94 $Y=1.557
+ $X2=6.195 $Y2=1.557
r88 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.94
+ $Y=1.515 $X2=5.94 $Y2=1.515
r89 45 47 22.1459 $w=3.7e-07 $l=1.7e-07 $layer=POLY_cond $X=5.77 $Y=1.557
+ $X2=5.94 $Y2=1.557
r90 44 45 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.745 $Y=1.557
+ $X2=5.77 $Y2=1.557
r91 43 44 52.7595 $w=3.7e-07 $l=4.05e-07 $layer=POLY_cond $X=5.34 $Y=1.557
+ $X2=5.745 $Y2=1.557
r92 42 43 5.86216 $w=3.7e-07 $l=4.5e-08 $layer=POLY_cond $X=5.295 $Y=1.557
+ $X2=5.34 $Y2=1.557
r93 40 42 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=4.92 $Y=1.557
+ $X2=5.295 $Y2=1.557
r94 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.92
+ $Y=1.515 $X2=4.92 $Y2=1.515
r95 38 40 1.3027 $w=3.7e-07 $l=1e-08 $layer=POLY_cond $X=4.91 $Y=1.557 $X2=4.92
+ $Y2=1.557
r96 37 38 8.46757 $w=3.7e-07 $l=6.5e-08 $layer=POLY_cond $X=4.845 $Y=1.557
+ $X2=4.91 $Y2=1.557
r97 32 48 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.94
+ $Y2=1.565
r98 31 48 11.2564 $w=4.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.94 $Y2=1.565
r99 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r100 30 41 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.92 $Y2=1.565
r101 29 41 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.92 $Y2=1.565
r102 25 50 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.2 $Y=1.35
+ $X2=6.2 $Y2=1.557
r103 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.2 $Y=1.35 $X2=6.2
+ $Y2=0.74
r104 22 49 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=1.557
r105 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=2.4
r106 18 45 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.77 $Y=1.35
+ $X2=5.77 $Y2=1.557
r107 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.77 $Y=1.35
+ $X2=5.77 $Y2=0.74
r108 15 44 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=1.557
r109 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=2.4
r110 11 43 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.34 $Y=1.35
+ $X2=5.34 $Y2=1.557
r111 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.34 $Y=1.35
+ $X2=5.34 $Y2=0.74
r112 8 42 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.295 $Y=1.765
+ $X2=5.295 $Y2=1.557
r113 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.295 $Y=1.765
+ $X2=5.295 $Y2=2.4
r114 4 38 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.91 $Y=1.35
+ $X2=4.91 $Y2=1.557
r115 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.91 $Y=1.35 $X2=4.91
+ $Y2=0.74
r116 1 37 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.845 $Y=1.765
+ $X2=4.845 $Y2=1.557
r117 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.845 $Y=1.765
+ $X2=4.845 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%B1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 47
c82 3 0 2.04552e-19 $X=6.63 $Y=0.74
r83 47 49 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=7.92 $Y=1.557
+ $X2=7.995 $Y2=1.557
r84 45 47 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=7.545 $Y=1.557
+ $X2=7.92 $Y2=1.557
r85 44 45 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=7.49 $Y=1.557
+ $X2=7.545 $Y2=1.557
r86 43 44 51.4568 $w=3.7e-07 $l=3.95e-07 $layer=POLY_cond $X=7.095 $Y=1.557
+ $X2=7.49 $Y2=1.557
r87 42 43 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=7.06 $Y=1.557
+ $X2=7.095 $Y2=1.557
r88 40 42 20.8432 $w=3.7e-07 $l=1.6e-07 $layer=POLY_cond $X=6.9 $Y=1.557
+ $X2=7.06 $Y2=1.557
r89 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.9
+ $Y=1.515 $X2=6.9 $Y2=1.515
r90 38 40 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=6.645 $Y=1.557
+ $X2=6.9 $Y2=1.557
r91 37 38 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=6.63 $Y=1.557
+ $X2=6.645 $Y2=1.557
r92 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.4 $Y2=1.565
r93 31 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.92
+ $Y=1.515 $X2=7.92 $Y2=1.515
r94 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r95 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r96 29 41 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=6.96 $Y=1.565 $X2=6.9
+ $Y2=1.565
r97 26 49 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.995 $Y=1.765
+ $X2=7.995 $Y2=1.557
r98 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.995 $Y=1.765
+ $X2=7.995 $Y2=2.4
r99 22 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.92 $Y=1.35
+ $X2=7.92 $Y2=1.557
r100 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.92 $Y=1.35
+ $X2=7.92 $Y2=0.74
r101 19 45 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.545 $Y=1.765
+ $X2=7.545 $Y2=1.557
r102 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.545 $Y=1.765
+ $X2=7.545 $Y2=2.4
r103 15 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.49 $Y=1.35
+ $X2=7.49 $Y2=1.557
r104 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.49 $Y=1.35
+ $X2=7.49 $Y2=0.74
r105 12 43 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.095 $Y=1.765
+ $X2=7.095 $Y2=1.557
r106 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.095 $Y=1.765
+ $X2=7.095 $Y2=2.4
r107 8 42 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.06 $Y=1.35
+ $X2=7.06 $Y2=1.557
r108 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.06 $Y=1.35
+ $X2=7.06 $Y2=0.74
r109 5 38 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.645 $Y=1.765
+ $X2=6.645 $Y2=1.557
r110 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.645 $Y=1.765
+ $X2=6.645 $Y2=2.4
r111 1 37 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=1.35
+ $X2=6.63 $Y2=1.557
r112 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.63 $Y=1.35 $X2=6.63
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%A_29_392# 1 2 3 12 16 17 18 21 22 24 26
r48 24 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.14 $X2=2.07
+ $Y2=2.055
r49 24 26 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.07 $Y=2.14
+ $X2=2.07 $Y2=2.815
r50 23 29 3.40825 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=1.255 $Y=2.055
+ $X2=1.17 $Y2=2.04
r51 22 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=2.055
+ $X2=2.07 $Y2=2.055
r52 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.905 $Y=2.055
+ $X2=1.255 $Y2=2.055
r53 19 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=2.905 $X2=1.17
+ $Y2=2.815
r54 18 29 3.40825 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.17 $Y=2.14 $X2=1.17
+ $Y2=2.04
r55 18 21 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.17 $Y=2.14
+ $X2=1.17 $Y2=2.815
r56 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.17 $Y2=2.905
r57 16 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.435 $Y2=2.99
r58 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.27 $Y=2.105
+ $X2=0.27 $Y2=2.815
r59 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.27 $Y=2.905
+ $X2=0.435 $Y2=2.99
r60 10 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=2.905 $X2=0.27
+ $Y2=2.815
r61 3 31 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.96 $X2=2.07 $Y2=2.135
r62 3 26 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.96 $X2=2.07 $Y2=2.815
r63 2 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.96 $X2=1.17 $Y2=2.105
r64 2 21 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.96 $X2=1.17 $Y2=2.815
r65 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.96 $X2=0.27 $Y2=2.815
r66 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.96 $X2=0.27 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%VPWR 1 2 3 4 5 18 20 24 28 32 36 39 40 42
+ 43 44 46 54 67 68 71 74 77
c106 18 0 1.88367e-19 $X=1.62 $Y=2.475
r107 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r108 74 75 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 71 72 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r111 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r112 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 62 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r115 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r116 59 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.01 $Y2=3.33
r117 59 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.48 $Y2=3.33
r118 58 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r119 58 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 55 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=3.33
+ $X2=5.07 $Y2=3.33
r122 55 57 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 54 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=6.01 $Y2=3.33
r124 54 57 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=5.52 $Y2=3.33
r125 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r126 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 49 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 48 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r129 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 46 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.455 $Y=3.33
+ $X2=1.58 $Y2=3.33
r131 46 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 44 75 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=5.04 $Y2=3.33
r133 44 72 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=1.68 $Y2=3.33
r134 42 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.685 $Y=3.33
+ $X2=7.44 $Y2=3.33
r135 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=3.33
+ $X2=7.77 $Y2=3.33
r136 41 67 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.855 $Y=3.33
+ $X2=8.4 $Y2=3.33
r137 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=3.33
+ $X2=7.77 $Y2=3.33
r138 39 61 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.48 $Y2=3.33
r139 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.83 $Y2=3.33
r140 38 64 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=7.44 $Y2=3.33
r141 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=6.83 $Y2=3.33
r142 34 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=3.245
+ $X2=7.77 $Y2=3.33
r143 34 36 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=7.77 $Y=3.245
+ $X2=7.77 $Y2=2.455
r144 30 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=3.33
r145 30 32 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=2.455
r146 26 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=3.33
r147 26 28 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.455
r148 22 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=3.245
+ $X2=5.07 $Y2=3.33
r149 22 24 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=5.07 $Y=3.245
+ $X2=5.07 $Y2=2.455
r150 21 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.58 $Y2=3.33
r151 20 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=5.07 $Y2=3.33
r152 20 21 213.989 $w=1.68e-07 $l=3.28e-06 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=1.705 $Y2=3.33
r153 16 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=3.245
+ $X2=1.58 $Y2=3.33
r154 16 18 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=1.58 $Y=3.245
+ $X2=1.58 $Y2=2.475
r155 5 36 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.62
+ $Y=1.84 $X2=7.77 $Y2=2.455
r156 4 32 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.72
+ $Y=1.84 $X2=6.87 $Y2=2.455
r157 3 28 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.82
+ $Y=1.84 $X2=5.97 $Y2=2.455
r158 2 24 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.92
+ $Y=1.84 $X2=5.07 $Y2=2.455
r159 1 18 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=1.96 $X2=1.62 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%A_539_368# 1 2 3 4 5 6 7 24 28 29 32 34 36
+ 39 40 44 46 50 52 56 58 60 62 64 68 70 72
c123 70 0 1.52151e-19 $X=6.42 $Y=1.985
r124 60 74 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.22 $Y=2.12 $X2=8.22
+ $Y2=2.035
r125 60 62 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.22 $Y=2.12
+ $X2=8.22 $Y2=2.815
r126 59 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=2.035
+ $X2=7.32 $Y2=2.035
r127 58 74 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.055 $Y=2.035
+ $X2=8.22 $Y2=2.035
r128 58 59 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.055 $Y=2.035
+ $X2=7.485 $Y2=2.035
r129 54 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.32 $Y=2.12
+ $X2=7.32 $Y2=2.035
r130 54 56 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.32 $Y=2.12
+ $X2=7.32 $Y2=2.815
r131 53 70 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=6.505 $Y=2.035
+ $X2=6.42 $Y2=1.97
r132 52 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.155 $Y=2.035
+ $X2=7.32 $Y2=2.035
r133 52 53 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.155 $Y=2.035
+ $X2=6.505 $Y2=2.035
r134 48 70 1.34256 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.42 $Y=2.12
+ $X2=6.42 $Y2=1.97
r135 48 50 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.42 $Y=2.12
+ $X2=6.42 $Y2=2.4
r136 47 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=2.035
+ $X2=5.52 $Y2=2.035
r137 46 70 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=6.335 $Y=2.035
+ $X2=6.42 $Y2=1.97
r138 46 47 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.335 $Y=2.035
+ $X2=5.685 $Y2=2.035
r139 42 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=2.12
+ $X2=5.52 $Y2=2.035
r140 42 44 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.52 $Y=2.12
+ $X2=5.52 $Y2=2.815
r141 41 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.785 $Y=2.035
+ $X2=4.62 $Y2=2.035
r142 40 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=2.035
+ $X2=5.52 $Y2=2.035
r143 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.355 $Y=2.035
+ $X2=4.785 $Y2=2.035
r144 37 39 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.62 $Y=2.905
+ $X2=4.62 $Y2=2.815
r145 36 66 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=2.12 $X2=4.62
+ $Y2=2.035
r146 36 39 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.62 $Y=2.12
+ $X2=4.62 $Y2=2.815
r147 35 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=2.99
+ $X2=3.72 $Y2=2.99
r148 34 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.455 $Y=2.99
+ $X2=4.62 $Y2=2.905
r149 34 35 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.455 $Y=2.99
+ $X2=3.885 $Y2=2.99
r150 30 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=2.905
+ $X2=3.72 $Y2=2.99
r151 30 32 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.72 $Y=2.905
+ $X2=3.72 $Y2=2.225
r152 28 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=2.99
+ $X2=3.72 $Y2=2.99
r153 28 29 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.555 $Y=2.99
+ $X2=2.985 $Y2=2.99
r154 24 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.82 $Y=1.985
+ $X2=2.82 $Y2=2.815
r155 22 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.82 $Y=2.905
+ $X2=2.985 $Y2=2.99
r156 22 27 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.82 $Y=2.905
+ $X2=2.82 $Y2=2.815
r157 7 74 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=1.84 $X2=8.22 $Y2=2.115
r158 7 62 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=1.84 $X2=8.22 $Y2=2.815
r159 6 72 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=7.17
+ $Y=1.84 $X2=7.32 $Y2=2.115
r160 6 56 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.17
+ $Y=1.84 $X2=7.32 $Y2=2.815
r161 5 70 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.84 $X2=6.42 $Y2=1.985
r162 5 50 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=6.27
+ $Y=1.84 $X2=6.42 $Y2=2.4
r163 4 68 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.37
+ $Y=1.84 $X2=5.52 $Y2=2.115
r164 4 44 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.37
+ $Y=1.84 $X2=5.52 $Y2=2.815
r165 3 66 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.84 $X2=4.62 $Y2=2.115
r166 3 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.84 $X2=4.62 $Y2=2.815
r167 2 32 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=3.57
+ $Y=1.84 $X2=3.72 $Y2=2.225
r168 1 27 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=1.84 $X2=2.82 $Y2=2.815
r169 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=1.84 $X2=2.82 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%Y 1 2 3 4 5 6 19 21 23 27 31 33 34 35 39
+ 43 45 50 52 55 56 57
c99 45 0 4.29123e-20 $X=5.985 $Y=0.95
c100 31 0 2.7959e-19 $X=3.295 $Y=0.515
c101 21 0 3.44467e-19 $X=2.435 $Y=0.515
c102 19 0 1.64164e-19 $X=2.395 $Y=0.79
r103 57 60 6.557 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=4.11 $Y=1.295
+ $X2=4.11 $Y2=1.13
r104 56 60 0.883768 $w=2.9e-07 $l=1.7e-07 $layer=LI1_cond $X=4.11 $Y=0.96
+ $X2=4.11 $Y2=1.13
r105 54 55 5.33064 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0.95
+ $X2=4.96 $Y2=0.95
r106 51 57 16.8893 $w=2.88e-07 $l=4.25e-07 $layer=LI1_cond $X=4.11 $Y=1.72
+ $X2=4.11 $Y2=1.295
r107 51 52 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=1.72
+ $X2=4.11 $Y2=1.805
r108 43 54 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=5.14 $Y=0.95
+ $X2=5.125 $Y2=0.95
r109 43 45 27.0504 $w=3.58e-07 $l=8.45e-07 $layer=LI1_cond $X=5.14 $Y=0.95
+ $X2=5.985 $Y2=0.95
r110 42 56 5.74179 $w=2.55e-07 $l=1.45e-07 $layer=LI1_cond $X=4.255 $Y=0.96
+ $X2=4.11 $Y2=0.96
r111 42 55 23.8962 $w=3.38e-07 $l=7.05e-07 $layer=LI1_cond $X=4.255 $Y=0.96
+ $X2=4.96 $Y2=0.96
r112 37 52 3.98977 $w=2.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.17 $Y=1.89
+ $X2=4.11 $Y2=1.805
r113 37 39 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.17 $Y=1.89
+ $X2=4.17 $Y2=1.985
r114 36 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.38 $Y=0.875
+ $X2=3.295 $Y2=0.875
r115 35 56 5.74179 $w=2.55e-07 $l=1.8262e-07 $layer=LI1_cond $X=3.965 $Y=0.875
+ $X2=4.11 $Y2=0.96
r116 35 36 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.965 $Y=0.875
+ $X2=3.38 $Y2=0.875
r117 33 52 2.45049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=4.11 $Y2=1.805
r118 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=3.355 $Y2=1.805
r119 29 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=0.79
+ $X2=3.295 $Y2=0.875
r120 29 31 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.295 $Y=0.79
+ $X2=3.295 $Y2=0.515
r121 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=1.89
+ $X2=3.355 $Y2=1.805
r122 25 27 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.27 $Y=1.89
+ $X2=3.27 $Y2=1.985
r123 24 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.52 $Y=0.875
+ $X2=2.395 $Y2=0.875
r124 23 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.875
+ $X2=3.295 $Y2=0.875
r125 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.21 $Y=0.875
+ $X2=2.52 $Y2=0.875
r126 19 48 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=0.79
+ $X2=2.395 $Y2=0.875
r127 19 21 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.395 $Y=0.79
+ $X2=2.395 $Y2=0.515
r128 6 39 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.02
+ $Y=1.84 $X2=4.17 $Y2=1.985
r129 5 27 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.12
+ $Y=1.84 $X2=3.27 $Y2=1.985
r130 4 45 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.37 $X2=5.985 $Y2=0.95
r131 3 54 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.985
+ $Y=0.37 $X2=5.125 $Y2=0.95
r132 2 50 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.37 $X2=3.295 $Y2=0.875
r133 2 31 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.37 $X2=3.295 $Y2=0.515
r134 1 48 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.37 $X2=2.435 $Y2=0.875
r135 1 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.37 $X2=2.435 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%VGND 1 2 3 4 5 6 21 25 29 31 35 39 43 46
+ 47 49 50 51 52 54 55 57 58 59 82 83 86
r111 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r112 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r113 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r114 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r115 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r116 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r117 74 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r118 73 76 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6.48
+ $Y2=0
r119 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r120 71 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.725
+ $Y2=0
r121 71 73 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.08
+ $Y2=0
r122 70 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r123 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r124 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r125 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r126 63 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r127 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r128 59 77 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=6.48 $Y2=0
r129 59 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r130 57 79 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=7.54 $Y=0 $X2=7.44
+ $Y2=0
r131 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.54 $Y=0 $X2=7.665
+ $Y2=0
r132 56 82 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.79 $Y=0 $X2=8.4
+ $Y2=0
r133 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.79 $Y=0 $X2=7.665
+ $Y2=0
r134 54 76 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.68 $Y=0 $X2=6.48
+ $Y2=0
r135 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.68 $Y=0 $X2=6.805
+ $Y2=0
r136 53 79 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.93 $Y=0 $X2=7.44
+ $Y2=0
r137 53 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.93 $Y=0 $X2=6.805
+ $Y2=0
r138 51 69 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.64
+ $Y2=0
r139 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.865
+ $Y2=0
r140 49 66 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=1.68
+ $Y2=0
r141 49 50 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=1.945
+ $Y2=0
r142 48 69 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.64
+ $Y2=0
r143 48 50 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.945
+ $Y2=0
r144 46 62 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=0.72
+ $Y2=0
r145 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=1.105
+ $Y2=0
r146 45 66 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.68
+ $Y2=0
r147 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.105
+ $Y2=0
r148 41 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=0.085
+ $X2=7.665 $Y2=0
r149 41 43 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=7.665 $Y=0.085
+ $X2=7.665 $Y2=0.675
r150 37 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=0.085
+ $X2=6.805 $Y2=0
r151 37 39 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=6.805 $Y=0.085
+ $X2=6.805 $Y2=0.675
r152 33 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0
r153 33 35 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0.525
r154 32 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.865
+ $Y2=0
r155 31 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=3.725
+ $Y2=0
r156 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=3.03
+ $Y2=0
r157 27 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0
r158 27 29 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0.525
r159 23 50 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=0.085
+ $X2=1.945 $Y2=0
r160 23 25 25.2345 $w=2.88e-07 $l=6.35e-07 $layer=LI1_cond $X=1.945 $Y=0.085
+ $X2=1.945 $Y2=0.72
r161 19 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=0.085
+ $X2=1.105 $Y2=0
r162 19 21 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.105 $Y=0.085
+ $X2=1.105 $Y2=0.525
r163 6 43 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=7.565
+ $Y=0.37 $X2=7.705 $Y2=0.675
r164 5 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.705
+ $Y=0.37 $X2=6.845 $Y2=0.675
r165 4 35 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.37 $X2=3.725 $Y2=0.525
r166 3 29 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.37 $X2=2.865 $Y2=0.525
r167 2 25 182 $w=1.7e-07 $l=4.22493e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.37 $X2=1.985 $Y2=0.72
r168 1 21 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.37 $X2=1.105 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_4%A_914_74# 1 2 3 4 5 16 22 26 27 30 32 36
+ 40
c54 26 0 1.52151e-19 $X=7.11 $Y=1.095
c55 22 0 1.6164e-19 $X=6.415 $Y=0.6
r56 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.135 $Y=1.01
+ $X2=8.135 $Y2=0.515
r57 33 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.36 $Y=1.095
+ $X2=7.235 $Y2=1.095
r58 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.97 $Y=1.095
+ $X2=8.135 $Y2=1.01
r59 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.97 $Y=1.095
+ $X2=7.36 $Y2=1.095
r60 28 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.235 $Y=1.01
+ $X2=7.235 $Y2=1.095
r61 28 30 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=7.235 $Y=1.01
+ $X2=7.235 $Y2=0.515
r62 26 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.11 $Y=1.095
+ $X2=7.235 $Y2=1.095
r63 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.11 $Y=1.095
+ $X2=6.5 $Y2=1.095
r64 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=1.01
+ $X2=6.5 $Y2=1.095
r65 23 25 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.415 $Y=1.01
+ $X2=6.415 $Y2=0.965
r66 22 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.415 $Y=0.6
+ $X2=6.415 $Y2=0.475
r67 22 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.415 $Y=0.6
+ $X2=6.415 $Y2=0.965
r68 18 21 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=4.695 $Y=0.475
+ $X2=5.555 $Y2=0.475
r69 16 39 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.33 $Y=0.475
+ $X2=6.415 $Y2=0.475
r70 16 21 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=6.33 $Y=0.475
+ $X2=5.555 $Y2=0.475
r71 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.995
+ $Y=0.37 $X2=8.135 $Y2=0.515
r72 4 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.135
+ $Y=0.37 $X2=7.275 $Y2=0.515
r73 3 39 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.275
+ $Y=0.37 $X2=6.415 $Y2=0.515
r74 3 25 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.275
+ $Y=0.37 $X2=6.415 $Y2=0.965
r75 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.37 $X2=5.555 $Y2=0.515
r76 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.37 $X2=4.695 $Y2=0.515
.ends

