* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__clkdlyinv3sd1_1 A VGND VNB VPB VPWR Y
M1000 VPWR A a_28_74# VPB pshort w=1.12e+06u l=150000u
+  ad=1.0448e+12p pd=6.44e+06u as=3.136e+11p ps=2.8e+06u
M1001 Y a_285_392# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1002 a_285_392# a_28_74# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1003 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=4.2e+11p pd=3.68e+06u as=1.113e+11p ps=1.37e+06u
M1004 a_285_392# a_28_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 Y a_285_392# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends
