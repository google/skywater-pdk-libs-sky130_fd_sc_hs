* File: sky130_fd_sc_hs__and3b_2.pxi.spice
* Created: Tue Sep  1 19:55:32 2020
* 
x_PM_SKY130_FD_SC_HS__AND3B_2%A_N N_A_N_c_76_n N_A_N_M1010_g N_A_N_c_81_n
+ N_A_N_M1008_g A_N N_A_N_c_78_n N_A_N_c_79_n PM_SKY130_FD_SC_HS__AND3B_2%A_N
x_PM_SKY130_FD_SC_HS__AND3B_2%A_27_88# N_A_27_88#_M1010_s N_A_27_88#_M1008_s
+ N_A_27_88#_c_107_n N_A_27_88#_c_115_n N_A_27_88#_M1005_g N_A_27_88#_c_108_n
+ N_A_27_88#_M1007_g N_A_27_88#_c_109_n N_A_27_88#_c_110_n N_A_27_88#_c_111_n
+ N_A_27_88#_c_112_n N_A_27_88#_c_117_n N_A_27_88#_c_113_n N_A_27_88#_c_114_n
+ N_A_27_88#_c_119_n N_A_27_88#_c_120_n N_A_27_88#_c_121_n
+ PM_SKY130_FD_SC_HS__AND3B_2%A_27_88#
x_PM_SKY130_FD_SC_HS__AND3B_2%B N_B_c_174_n N_B_M1006_g N_B_c_175_n N_B_M1003_g
+ B B B B PM_SKY130_FD_SC_HS__AND3B_2%B
x_PM_SKY130_FD_SC_HS__AND3B_2%C N_C_M1000_g N_C_c_211_n N_C_M1004_g C
+ PM_SKY130_FD_SC_HS__AND3B_2%C
x_PM_SKY130_FD_SC_HS__AND3B_2%A_284_368# N_A_284_368#_M1007_s
+ N_A_284_368#_M1005_s N_A_284_368#_M1003_d N_A_284_368#_M1002_g
+ N_A_284_368#_c_249_n N_A_284_368#_M1001_g N_A_284_368#_M1011_g
+ N_A_284_368#_c_250_n N_A_284_368#_M1009_g N_A_284_368#_c_245_n
+ N_A_284_368#_c_252_n N_A_284_368#_c_268_n N_A_284_368#_c_253_n
+ N_A_284_368#_c_254_n N_A_284_368#_c_246_n N_A_284_368#_c_256_n
+ N_A_284_368#_c_272_n N_A_284_368#_c_247_n N_A_284_368#_c_248_n
+ PM_SKY130_FD_SC_HS__AND3B_2%A_284_368#
x_PM_SKY130_FD_SC_HS__AND3B_2%VPWR N_VPWR_M1008_d N_VPWR_M1005_d N_VPWR_M1004_d
+ N_VPWR_M1009_d N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n
+ N_VPWR_c_348_n N_VPWR_c_349_n N_VPWR_c_350_n VPWR N_VPWR_c_351_n
+ N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_343_n
+ PM_SKY130_FD_SC_HS__AND3B_2%VPWR
x_PM_SKY130_FD_SC_HS__AND3B_2%X N_X_M1002_d N_X_M1001_s N_X_c_399_n X X X X X
+ PM_SKY130_FD_SC_HS__AND3B_2%X
x_PM_SKY130_FD_SC_HS__AND3B_2%VGND N_VGND_M1010_d N_VGND_M1000_d N_VGND_M1011_s
+ N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n N_VGND_c_431_n
+ N_VGND_c_432_n VGND N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n
+ N_VGND_c_436_n PM_SKY130_FD_SC_HS__AND3B_2%VGND
cc_1 VNB N_A_N_c_76_n 0.0195074f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.755
cc_2 VNB N_A_N_M1010_g 0.0372275f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.715
cc_3 VNB N_A_N_c_78_n 0.0204063f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.425
cc_4 VNB N_A_N_c_79_n 0.0162384f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.425
cc_5 VNB N_A_27_88#_c_107_n 0.0559453f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_6 VNB N_A_27_88#_c_108_n 0.0196408f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.425
cc_7 VNB N_A_27_88#_c_109_n 0.0200972f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.26
cc_8 VNB N_A_27_88#_c_110_n 0.0211815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_88#_c_111_n 0.0283998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_88#_c_112_n 0.00959922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_88#_c_113_n 0.00179898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_88#_c_114_n 0.0375386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_174_n 0.0174585f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.435
cc_14 VNB N_B_c_175_n 0.0366156f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.715
cc_15 VNB B 0.00518004f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_16 VNB N_C_M1000_g 0.0266942f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.26
cc_17 VNB N_C_c_211_n 0.0226109f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.715
cc_18 VNB C 0.00914442f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_19 VNB N_A_284_368#_M1002_g 0.0230215f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.425
cc_20 VNB N_A_284_368#_M1011_g 0.0260225f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.595
cc_21 VNB N_A_284_368#_c_245_n 0.0191617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_284_368#_c_246_n 0.00121168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_284_368#_c_247_n 0.00753363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_284_368#_c_248_n 0.0928541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_343_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.425
cc_27 VNB X 0.00185591f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.425
cc_28 VNB N_VGND_c_427_n 0.0185992f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.425
cc_29 VNB N_VGND_c_428_n 0.00925448f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.595
cc_30 VNB N_VGND_c_429_n 0.0125919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_430_n 0.0419252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_431_n 0.0561173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_432_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_433_n 0.0177296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_434_n 0.0212406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_435_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_436_n 0.289569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_N_c_76_n 0.040174f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.755
cc_39 VPB N_A_N_c_81_n 0.0224362f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_40 VPB N_A_N_c_79_n 0.0112383f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.425
cc_41 VPB N_A_27_88#_c_115_n 0.0194225f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_42 VPB N_A_27_88#_c_109_n 0.00725985f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.26
cc_43 VPB N_A_27_88#_c_117_n 0.0211132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_27_88#_c_114_n 0.0249773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_27_88#_c_119_n 0.0051971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_27_88#_c_120_n 0.0386723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_88#_c_121_n 0.00647567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_B_c_175_n 0.0225969f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.715
cc_49 VPB B 0.00343199f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_50 VPB N_C_c_211_n 0.0262717f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.715
cc_51 VPB C 0.00707012f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_52 VPB N_A_284_368#_c_249_n 0.017011f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.425
cc_53 VPB N_A_284_368#_c_250_n 0.0172687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_284_368#_c_245_n 0.00257159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_284_368#_c_252_n 0.0181936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_284_368#_c_253_n 0.003137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_284_368#_c_254_n 0.00769764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_284_368#_c_246_n 0.0218388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_284_368#_c_256_n 0.00217379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_284_368#_c_248_n 0.0135395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_344_n 0.0204506f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.26
cc_62 VPB N_VPWR_c_345_n 0.0198956f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.595
cc_63 VPB N_VPWR_c_346_n 0.0103692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_347_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_348_n 0.0240489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_349_n 0.0297343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_350_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_351_n 0.017913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_352_n 0.0211424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_353_n 0.0182362f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_354_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_355_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_343_n 0.102248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_X_c_399_n 2.45031e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_75 VPB X 0.00115925f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.425
cc_76 N_A_N_M1010_g N_A_27_88#_c_110_n 0.00218986f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_77 N_A_N_M1010_g N_A_27_88#_c_111_n 0.0180286f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_78 N_A_N_c_78_n N_A_27_88#_c_111_n 0.00116829f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_79 N_A_N_c_79_n N_A_27_88#_c_111_n 0.0133787f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_80 N_A_N_c_78_n N_A_27_88#_c_112_n 0.00415347f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_81 N_A_N_c_79_n N_A_27_88#_c_112_n 0.022566f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_82 N_A_N_c_76_n N_A_27_88#_c_117_n 8.39929e-19 $X=0.395 $Y=1.755 $X2=0 $Y2=0
cc_83 N_A_N_c_81_n N_A_27_88#_c_117_n 0.0157224f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_84 N_A_N_c_79_n N_A_27_88#_c_117_n 0.0114298f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_85 N_A_N_M1010_g N_A_27_88#_c_113_n 0.00441126f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_86 N_A_N_c_79_n N_A_27_88#_c_113_n 0.0287652f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_87 N_A_N_M1010_g N_A_27_88#_c_114_n 0.0250202f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_88 N_A_N_c_79_n N_A_27_88#_c_114_n 0.00256857f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_89 N_A_N_c_76_n N_A_27_88#_c_119_n 0.00650482f $X=0.395 $Y=1.755 $X2=0 $Y2=0
cc_90 N_A_N_c_76_n N_A_27_88#_c_120_n 0.00483226f $X=0.395 $Y=1.755 $X2=0 $Y2=0
cc_91 N_A_N_c_81_n N_A_27_88#_c_120_n 0.003607f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_92 N_A_N_c_79_n N_A_27_88#_c_120_n 0.0248079f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_93 N_A_N_c_78_n N_A_27_88#_c_121_n 0.00145659f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_94 N_A_N_c_81_n N_VPWR_c_344_n 0.0159649f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_95 N_A_N_c_81_n N_VPWR_c_351_n 0.00429299f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_96 N_A_N_c_81_n N_VPWR_c_343_n 0.00851215f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_97 N_A_N_M1010_g N_VGND_c_427_n 0.0117471f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_98 N_A_N_M1010_g N_VGND_c_433_n 0.00438299f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_99 N_A_N_M1010_g N_VGND_c_436_n 0.00439883f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_100 N_A_27_88#_c_108_n N_B_c_174_n 0.0342483f $X=1.805 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_27_88#_c_115_n N_B_c_175_n 0.0269757f $X=1.79 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_27_88#_c_109_n N_B_c_175_n 0.0399506f $X=1.79 $Y=1.475 $X2=0 $Y2=0
cc_103 N_A_27_88#_c_108_n B 0.0106431f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_104 N_A_27_88#_c_107_n N_A_284_368#_c_245_n 0.0327021f $X=1.7 $Y=1.397 $X2=0
+ $Y2=0
cc_105 N_A_27_88#_c_115_n N_A_284_368#_c_245_n 0.00491791f $X=1.79 $Y=1.765
+ $X2=0 $Y2=0
cc_106 N_A_27_88#_c_108_n N_A_284_368#_c_245_n 0.0144396f $X=1.805 $Y=1.185
+ $X2=0 $Y2=0
cc_107 N_A_27_88#_c_109_n N_A_284_368#_c_245_n 0.012456f $X=1.79 $Y=1.475 $X2=0
+ $Y2=0
cc_108 N_A_27_88#_c_111_n N_A_284_368#_c_245_n 0.0151173f $X=0.9 $Y=1.005 $X2=0
+ $Y2=0
cc_109 N_A_27_88#_c_113_n N_A_284_368#_c_245_n 0.059451f $X=1.065 $Y=1.35 $X2=0
+ $Y2=0
cc_110 N_A_27_88#_c_114_n N_A_284_368#_c_245_n 0.00218282f $X=1.065 $Y=1.35
+ $X2=0 $Y2=0
cc_111 N_A_27_88#_c_119_n N_A_284_368#_c_245_n 0.00473674f $X=0.985 $Y=2.1 $X2=0
+ $Y2=0
cc_112 N_A_27_88#_c_115_n N_A_284_368#_c_252_n 0.00937054f $X=1.79 $Y=1.765
+ $X2=0 $Y2=0
cc_113 N_A_27_88#_c_117_n N_A_284_368#_c_252_n 0.00834063f $X=0.9 $Y=2.185 $X2=0
+ $Y2=0
cc_114 N_A_27_88#_c_115_n N_A_284_368#_c_268_n 0.0140213f $X=1.79 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_27_88#_c_115_n N_A_284_368#_c_256_n 0.00187028f $X=1.79 $Y=1.765
+ $X2=0 $Y2=0
cc_116 N_A_27_88#_c_117_n N_A_284_368#_c_256_n 0.00117914f $X=0.9 $Y=2.185 $X2=0
+ $Y2=0
cc_117 N_A_27_88#_c_119_n N_A_284_368#_c_256_n 0.00796474f $X=0.985 $Y=2.1 $X2=0
+ $Y2=0
cc_118 N_A_27_88#_c_115_n N_A_284_368#_c_272_n 9.66317e-19 $X=1.79 $Y=1.765
+ $X2=0 $Y2=0
cc_119 N_A_27_88#_c_117_n N_VPWR_M1008_d 0.00366719f $X=0.9 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_27_88#_c_117_n N_VPWR_c_344_n 0.0220028f $X=0.9 $Y=2.185 $X2=0 $Y2=0
cc_121 N_A_27_88#_c_120_n N_VPWR_c_344_n 0.0210352f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_122 N_A_27_88#_c_115_n N_VPWR_c_345_n 0.00685345f $X=1.79 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_27_88#_c_115_n N_VPWR_c_349_n 0.00481995f $X=1.79 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_27_88#_c_120_n N_VPWR_c_351_n 0.0126277f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_125 N_A_27_88#_c_115_n N_VPWR_c_343_n 0.00508379f $X=1.79 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_27_88#_c_120_n N_VPWR_c_343_n 0.0104521f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_127 N_A_27_88#_c_111_n N_VGND_M1010_d 0.00296919f $X=0.9 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_27_88#_c_110_n N_VGND_c_427_n 0.0131449f $X=0.28 $Y=0.715 $X2=0 $Y2=0
cc_129 N_A_27_88#_c_111_n N_VGND_c_427_n 0.0219096f $X=0.9 $Y=1.005 $X2=0 $Y2=0
cc_130 N_A_27_88#_c_108_n N_VGND_c_431_n 0.00434272f $X=1.805 $Y=1.185 $X2=0
+ $Y2=0
cc_131 N_A_27_88#_c_110_n N_VGND_c_433_n 0.0089644f $X=0.28 $Y=0.715 $X2=0 $Y2=0
cc_132 N_A_27_88#_c_108_n N_VGND_c_436_n 0.00825979f $X=1.805 $Y=1.185 $X2=0
+ $Y2=0
cc_133 N_A_27_88#_c_110_n N_VGND_c_436_n 0.00911107f $X=0.28 $Y=0.715 $X2=0
+ $Y2=0
cc_134 N_B_c_174_n N_C_M1000_g 0.0240719f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_135 N_B_c_175_n N_C_M1000_g 0.0245655f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_136 B N_C_M1000_g 0.00907035f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_137 N_B_c_175_n N_C_c_211_n 0.012263f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_138 B N_C_c_211_n 5.73912e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_139 N_B_c_175_n C 0.0017578f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_140 B C 0.0263467f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_141 N_B_c_174_n N_A_284_368#_c_245_n 0.00150231f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_142 N_B_c_175_n N_A_284_368#_c_245_n 9.78495e-19 $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_143 B N_A_284_368#_c_245_n 0.0716531f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_144 N_B_c_175_n N_A_284_368#_c_252_n 8.71718e-19 $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_145 N_B_c_175_n N_A_284_368#_c_268_n 0.0136588f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_146 B N_A_284_368#_c_268_n 0.0280724f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_147 N_B_c_175_n N_A_284_368#_c_253_n 0.00495314f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_148 N_B_c_175_n N_A_284_368#_c_272_n 0.0054806f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_149 B N_A_284_368#_c_272_n 0.00179867f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_150 N_B_c_175_n N_VPWR_c_345_n 0.00663439f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_151 N_B_c_175_n N_VPWR_c_352_n 0.00481995f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_152 N_B_c_175_n N_VPWR_c_343_n 0.00508379f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_153 N_B_c_174_n N_VGND_c_428_n 0.0015178f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_154 B N_VGND_c_428_n 0.030309f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_155 N_B_c_174_n N_VGND_c_431_n 0.00303293f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_156 B N_VGND_c_431_n 0.0108342f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_157 N_B_c_174_n N_VGND_c_436_n 0.00372643f $X=2.195 $Y=1.22 $X2=0 $Y2=0
cc_158 B N_VGND_c_436_n 0.0133038f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_159 B A_376_74# 0.00738039f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_160 B A_454_74# 0.00983395f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_161 N_C_M1000_g N_A_284_368#_M1002_g 0.0181973f $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_162 N_C_c_211_n N_A_284_368#_c_249_n 0.029368f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_163 N_C_c_211_n N_A_284_368#_c_253_n 0.00660631f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_164 N_C_c_211_n N_A_284_368#_c_254_n 0.0145072f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_165 C N_A_284_368#_c_254_n 0.0168221f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_166 N_C_c_211_n N_A_284_368#_c_272_n 0.00651386f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_167 C N_A_284_368#_c_272_n 0.00305544f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_168 N_C_c_211_n N_A_284_368#_c_248_n 0.0203031f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_169 C N_A_284_368#_c_248_n 0.00390334f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_170 N_C_c_211_n N_VPWR_c_346_n 0.00561364f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_171 N_C_c_211_n N_VPWR_c_352_n 0.00481995f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_172 N_C_c_211_n N_VPWR_c_343_n 0.00508379f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_173 N_C_M1000_g X 2.59942e-19 $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_174 N_C_M1000_g X 2.16826e-19 $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_175 N_C_c_211_n X 0.00144181f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_176 C X 0.034443f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_177 N_C_M1000_g N_VGND_c_428_n 0.0179953f $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_178 N_C_c_211_n N_VGND_c_428_n 0.00426817f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_179 C N_VGND_c_428_n 0.0236581f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_180 N_C_M1000_g N_VGND_c_431_n 0.00383152f $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_181 N_C_M1000_g N_VGND_c_436_n 0.00758792f $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_284_368#_c_268_n N_VPWR_M1005_d 0.0103145f $X=2.42 $Y=2.035 $X2=0
+ $Y2=0
cc_183 N_A_284_368#_c_254_n N_VPWR_M1004_d 0.00832612f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_184 N_A_284_368#_c_254_n N_VPWR_M1009_d 0.00523446f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_185 N_A_284_368#_c_246_n N_VPWR_M1009_d 0.00715176f $X=4.13 $Y=2.24 $X2=0
+ $Y2=0
cc_186 N_A_284_368#_c_252_n N_VPWR_c_344_n 0.0165803f $X=1.565 $Y=2.695 $X2=0
+ $Y2=0
cc_187 N_A_284_368#_c_252_n N_VPWR_c_345_n 0.0221782f $X=1.565 $Y=2.695 $X2=0
+ $Y2=0
cc_188 N_A_284_368#_c_268_n N_VPWR_c_345_n 0.0248957f $X=2.42 $Y=2.035 $X2=0
+ $Y2=0
cc_189 N_A_284_368#_c_272_n N_VPWR_c_345_n 0.020261f $X=2.585 $Y=2.035 $X2=0
+ $Y2=0
cc_190 N_A_284_368#_c_249_n N_VPWR_c_346_n 0.0127815f $X=3.35 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A_284_368#_c_250_n N_VPWR_c_346_n 0.00152188f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_284_368#_c_253_n N_VPWR_c_346_n 0.0185061f $X=2.585 $Y=2.715 $X2=0
+ $Y2=0
cc_193 N_A_284_368#_c_254_n N_VPWR_c_346_n 0.0219335f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_194 N_A_284_368#_c_249_n N_VPWR_c_348_n 0.00152188f $X=3.35 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_284_368#_c_250_n N_VPWR_c_348_n 0.0132257f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_284_368#_c_254_n N_VPWR_c_348_n 0.0233188f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_197 N_A_284_368#_c_252_n N_VPWR_c_349_n 0.0097982f $X=1.565 $Y=2.695 $X2=0
+ $Y2=0
cc_198 N_A_284_368#_c_253_n N_VPWR_c_352_n 0.00976219f $X=2.585 $Y=2.715 $X2=0
+ $Y2=0
cc_199 N_A_284_368#_c_249_n N_VPWR_c_353_n 0.00413917f $X=3.35 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_284_368#_c_250_n N_VPWR_c_353_n 0.00413917f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A_284_368#_c_249_n N_VPWR_c_343_n 0.00817869f $X=3.35 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_284_368#_c_250_n N_VPWR_c_343_n 0.00817869f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_284_368#_c_252_n N_VPWR_c_343_n 0.0111907f $X=1.565 $Y=2.695 $X2=0
+ $Y2=0
cc_204 N_A_284_368#_c_253_n N_VPWR_c_343_n 0.0111764f $X=2.585 $Y=2.715 $X2=0
+ $Y2=0
cc_205 N_A_284_368#_c_254_n N_X_M1001_s 0.00962813f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_206 N_A_284_368#_c_249_n N_X_c_399_n 0.00526973f $X=3.35 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A_284_368#_c_250_n N_X_c_399_n 0.00435114f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_284_368#_c_254_n N_X_c_399_n 0.0183244f $X=4.045 $Y=2.325 $X2=0 $Y2=0
cc_209 N_A_284_368#_c_246_n N_X_c_399_n 0.0123189f $X=4.13 $Y=2.24 $X2=0 $Y2=0
cc_210 N_A_284_368#_c_272_n N_X_c_399_n 0.00291129f $X=2.585 $Y=2.035 $X2=0
+ $Y2=0
cc_211 N_A_284_368#_c_248_n N_X_c_399_n 0.00115735f $X=3.815 $Y=1.532 $X2=0
+ $Y2=0
cc_212 N_A_284_368#_M1002_g X 0.00855013f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_284_368#_M1011_g X 0.00788704f $X=3.765 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_284_368#_M1002_g X 0.00345332f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_284_368#_M1011_g X 0.00202916f $X=3.765 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_284_368#_M1002_g X 0.00483694f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_284_368#_c_249_n X 0.00147523f $X=3.35 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_284_368#_M1011_g X 0.00892301f $X=3.765 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_284_368#_c_250_n X 5.97294e-19 $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_284_368#_c_246_n X 0.00937974f $X=4.13 $Y=2.24 $X2=0 $Y2=0
cc_221 N_A_284_368#_c_247_n X 0.0246163f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_222 N_A_284_368#_c_248_n X 0.0305635f $X=3.815 $Y=1.532 $X2=0 $Y2=0
cc_223 N_A_284_368#_c_245_n N_VGND_c_427_n 0.0153399f $X=1.59 $Y=0.515 $X2=0
+ $Y2=0
cc_224 N_A_284_368#_M1002_g N_VGND_c_428_n 0.0100794f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_284_368#_M1011_g N_VGND_c_430_n 0.00647412f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_A_284_368#_c_247_n N_VGND_c_430_n 0.0214533f $X=4.05 $Y=1.465 $X2=0
+ $Y2=0
cc_227 N_A_284_368#_c_248_n N_VGND_c_430_n 0.00196248f $X=3.815 $Y=1.532 $X2=0
+ $Y2=0
cc_228 N_A_284_368#_c_245_n N_VGND_c_431_n 0.0156794f $X=1.59 $Y=0.515 $X2=0
+ $Y2=0
cc_229 N_A_284_368#_M1002_g N_VGND_c_434_n 0.00434272f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_230 N_A_284_368#_M1011_g N_VGND_c_434_n 0.00434272f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_231 N_A_284_368#_M1002_g N_VGND_c_436_n 0.00822522f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_284_368#_M1011_g N_VGND_c_436_n 0.0082413f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_284_368#_c_245_n N_VGND_c_436_n 0.0129217f $X=1.59 $Y=0.515 $X2=0
+ $Y2=0
cc_234 X N_VGND_c_428_n 0.0465051f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_235 X N_VGND_c_430_n 0.0293763f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_236 X N_VGND_c_434_n 0.0144922f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_237 X N_VGND_c_436_n 0.0118826f $X=3.515 $Y=0.47 $X2=0 $Y2=0
