* File: sky130_fd_sc_hs__clkinv_2.spice
* Created: Thu Aug 27 20:37:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__clkinv_2.pex.spice"
.subckt sky130_fd_sc_hs__clkinv_2  VNB VPB A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.1638 PD=1.41 PS=1.2 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.1638 PD=1.41 PS=1.2 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.3304
+ AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75001.1 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1003_d N_A_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.1
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX5_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_hs__clkinv_2.pxi.spice"
*
.ends
*
*
