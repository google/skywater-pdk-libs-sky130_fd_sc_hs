* File: sky130_fd_sc_hs__and3b_4.pxi.spice
* Created: Thu Aug 27 20:32:55 2020
* 
x_PM_SKY130_FD_SC_HS__AND3B_4%A_N N_A_N_M1020_g N_A_N_c_125_n N_A_N_M1010_g A_N
+ PM_SKY130_FD_SC_HS__AND3B_4%A_N
x_PM_SKY130_FD_SC_HS__AND3B_4%A_27_74# N_A_27_74#_M1020_s N_A_27_74#_M1010_s
+ N_A_27_74#_c_162_n N_A_27_74#_M1004_g N_A_27_74#_M1000_g N_A_27_74#_c_163_n
+ N_A_27_74#_M1008_g N_A_27_74#_M1018_g N_A_27_74#_c_157_n N_A_27_74#_c_158_n
+ N_A_27_74#_c_165_n N_A_27_74#_c_166_n N_A_27_74#_c_167_n N_A_27_74#_c_168_n
+ N_A_27_74#_c_159_n N_A_27_74#_c_169_n N_A_27_74#_c_160_n N_A_27_74#_c_161_n
+ PM_SKY130_FD_SC_HS__AND3B_4%A_27_74#
x_PM_SKY130_FD_SC_HS__AND3B_4%B N_B_M1015_g N_B_c_245_n N_B_M1001_g N_B_c_246_n
+ N_B_M1007_g N_B_M1016_g B B N_B_c_244_n PM_SKY130_FD_SC_HS__AND3B_4%B
x_PM_SKY130_FD_SC_HS__AND3B_4%C N_C_c_302_n N_C_M1019_g N_C_c_297_n N_C_M1003_g
+ N_C_c_303_n N_C_M1021_g N_C_c_298_n N_C_c_299_n N_C_c_300_n N_C_M1014_g C
+ N_C_c_301_n PM_SKY130_FD_SC_HS__AND3B_4%C
x_PM_SKY130_FD_SC_HS__AND3B_4%A_298_368# N_A_298_368#_M1000_s
+ N_A_298_368#_M1004_d N_A_298_368#_M1001_d N_A_298_368#_M1019_d
+ N_A_298_368#_c_366_n N_A_298_368#_M1002_g N_A_298_368#_c_355_n
+ N_A_298_368#_c_356_n N_A_298_368#_M1006_g N_A_298_368#_c_369_n
+ N_A_298_368#_M1005_g N_A_298_368#_M1011_g N_A_298_368#_c_370_n
+ N_A_298_368#_M1009_g N_A_298_368#_M1013_g N_A_298_368#_c_371_n
+ N_A_298_368#_M1012_g N_A_298_368#_M1017_g N_A_298_368#_c_372_n
+ N_A_298_368#_c_527_p N_A_298_368#_c_382_n N_A_298_368#_c_373_n
+ N_A_298_368#_c_402_n N_A_298_368#_c_374_n N_A_298_368#_c_375_n
+ N_A_298_368#_c_424_n N_A_298_368#_c_361_n N_A_298_368#_c_484_p
+ N_A_298_368#_c_376_n N_A_298_368#_c_362_n N_A_298_368#_c_363_n
+ N_A_298_368#_c_407_n N_A_298_368#_c_427_n N_A_298_368#_c_364_n
+ N_A_298_368#_c_365_n PM_SKY130_FD_SC_HS__AND3B_4%A_298_368#
x_PM_SKY130_FD_SC_HS__AND3B_4%VPWR N_VPWR_M1010_d N_VPWR_M1008_s N_VPWR_M1007_s
+ N_VPWR_M1021_s N_VPWR_M1005_s N_VPWR_M1012_s N_VPWR_c_534_n N_VPWR_c_535_n
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n
+ N_VPWR_c_541_n N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n VPWR
+ N_VPWR_c_545_n N_VPWR_c_546_n N_VPWR_c_547_n N_VPWR_c_548_n N_VPWR_c_533_n
+ N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n N_VPWR_c_553_n
+ PM_SKY130_FD_SC_HS__AND3B_4%VPWR
x_PM_SKY130_FD_SC_HS__AND3B_4%X N_X_M1006_s N_X_M1013_s N_X_M1002_d N_X_M1009_d
+ N_X_c_638_n N_X_c_639_n N_X_c_640_n N_X_c_631_n N_X_c_632_n N_X_c_633_n
+ N_X_c_641_n N_X_c_634_n N_X_c_635_n N_X_c_643_n N_X_c_644_n N_X_c_636_n X
+ PM_SKY130_FD_SC_HS__AND3B_4%X
x_PM_SKY130_FD_SC_HS__AND3B_4%VGND N_VGND_M1020_d N_VGND_M1003_s N_VGND_M1014_s
+ N_VGND_M1011_d N_VGND_M1017_d N_VGND_c_716_n N_VGND_c_717_n N_VGND_c_718_n
+ N_VGND_c_719_n N_VGND_c_720_n N_VGND_c_721_n VGND N_VGND_c_722_n
+ N_VGND_c_723_n N_VGND_c_724_n N_VGND_c_725_n N_VGND_c_726_n N_VGND_c_727_n
+ N_VGND_c_728_n N_VGND_c_729_n N_VGND_c_730_n N_VGND_c_731_n
+ PM_SKY130_FD_SC_HS__AND3B_4%VGND
x_PM_SKY130_FD_SC_HS__AND3B_4%A_239_98# N_A_239_98#_M1000_d N_A_239_98#_M1018_d
+ N_A_239_98#_M1016_d N_A_239_98#_c_808_n N_A_239_98#_c_809_n
+ N_A_239_98#_c_810_n N_A_239_98#_c_811_n N_A_239_98#_c_812_n
+ N_A_239_98#_c_813_n PM_SKY130_FD_SC_HS__AND3B_4%A_239_98#
x_PM_SKY130_FD_SC_HS__AND3B_4%A_498_98# N_A_498_98#_M1015_s N_A_498_98#_M1003_d
+ N_A_498_98#_c_853_n N_A_498_98#_c_854_n N_A_498_98#_c_855_n
+ PM_SKY130_FD_SC_HS__AND3B_4%A_498_98#
cc_1 VNB N_A_N_M1020_g 0.0276194f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_A_N_c_125_n 0.0663309f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.765
cc_3 VNB A_N 0.0062237f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_27_74#_M1000_g 0.0240643f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.345
cc_5 VNB N_A_27_74#_M1018_g 0.0197626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_74#_c_157_n 0.0214427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_c_158_n 0.0316559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_159_n 0.00745004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_160_n 0.00847386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_161_n 0.0650323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_M1015_g 0.0224581f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_12 VNB N_B_M1016_g 0.0253169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB B 0.00380401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_c_244_n 0.0373495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C_c_297_n 0.0181081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C_c_298_n 0.0213458f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.345
cc_17 VNB N_C_c_299_n 0.0699208f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.345
cc_18 VNB N_C_c_300_n 0.0160701f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.345
cc_19 VNB N_C_c_301_n 0.00465705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_298_368#_c_355_n 0.00543726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_298_368#_c_356_n 0.00772026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_298_368#_M1006_g 0.0237886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_298_368#_M1011_g 0.0214712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_298_368#_M1013_g 0.0205514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_298_368#_M1017_g 0.0276849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_298_368#_c_361_n 0.00498716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_298_368#_c_362_n 0.00316361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_298_368#_c_363_n 4.21191e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_298_368#_c_364_n 0.0144156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_298_368#_c_365_n 0.0933497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_533_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_631_n 0.00252795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_632_n 0.00369082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_633_n 0.00195434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_634_n 0.00187814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_635_n 0.0074247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_636_n 2.809e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB X 0.00857289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_716_n 0.017312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_717_n 0.017155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_718_n 0.00942615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_719_n 0.00262969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_720_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_721_n 0.0428762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_722_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_723_n 0.0673449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_724_n 0.0177559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_725_n 0.0167762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_726_n 0.0157319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_727_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_728_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_729_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_730_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_731_n 0.396591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_239_98#_c_808_n 0.0102458f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.345
cc_56 VNB N_A_239_98#_c_809_n 0.00919954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_239_98#_c_810_n 0.00478547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_239_98#_c_811_n 0.00919485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_239_98#_c_812_n 0.00659787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_239_98#_c_813_n 0.00273295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_498_98#_c_853_n 0.0197357f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=2.34
cc_62 VNB N_A_498_98#_c_854_n 0.00241395f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.345
cc_63 VNB N_A_498_98#_c_855_n 0.00517884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_A_N_c_125_n 0.0271957f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.765
cc_65 VPB N_A_27_74#_c_162_n 0.0155995f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=2.34
cc_66 VPB N_A_27_74#_c_163_n 0.0154109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_74#_c_158_n 0.00101234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_27_74#_c_165_n 0.0101156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_74#_c_166_n 0.0148348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_74#_c_167_n 0.0416815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_74#_c_168_n 0.00614929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_74#_c_169_n 0.00267435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_74#_c_160_n 0.00162357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_27_74#_c_161_n 0.0137268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_B_c_245_n 0.015627f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.765
cc_76 VPB N_B_c_246_n 0.0161028f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_77 VPB B 0.00702457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_B_c_244_n 0.0206013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_C_c_302_n 0.0159797f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.18
cc_80 VPB N_C_c_303_n 0.0156309f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=2.34
cc_81 VPB N_C_c_299_n 0.0256915f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.345
cc_82 VPB N_C_c_301_n 0.0048502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_298_368#_c_366_n 0.0164086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_298_368#_c_355_n 0.00463449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_298_368#_c_356_n 0.0059473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_298_368#_c_369_n 0.0159605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_298_368#_c_370_n 0.0159564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_298_368#_c_371_n 0.0166102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_298_368#_c_372_n 0.003137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_298_368#_c_373_n 0.003137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_298_368#_c_374_n 0.003137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_298_368#_c_375_n 0.00118251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_298_368#_c_376_n 0.00211648f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_298_368#_c_362_n 0.00129032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_298_368#_c_365_n 0.0385915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_534_n 0.0165851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_535_n 0.0133429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_536_n 0.0166833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_537_n 0.0220402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_538_n 0.0163399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_539_n 0.00830446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_540_n 0.0438947f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_541_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_542_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_543_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_544_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_545_n 0.0311457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_546_n 0.0192331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_547_n 0.0192331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_548_n 0.0123263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_533_n 0.121745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_550_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_551_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_552_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_553_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_X_c_638_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_X_c_639_n 0.00236064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_X_c_640_n 0.0017746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_X_c_641_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_X_c_635_n 0.0011613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_X_c_643_n 0.00355938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_X_c_644_n 0.00209569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB X 0.0221609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 N_A_N_c_125_n N_A_27_74#_c_162_n 0.0259731f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_N_c_125_n N_A_27_74#_M1000_g 0.00351198f $X=0.865 $Y=1.765 $X2=0
+ $Y2=0
cc_126 A_N N_A_27_74#_M1000_g 6.2207e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A_N_M1020_g N_A_27_74#_c_157_n 0.00588436f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_128 N_A_N_M1020_g N_A_27_74#_c_158_n 0.0146145f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_129 N_A_N_c_125_n N_A_27_74#_c_158_n 0.00423463f $X=0.865 $Y=1.765 $X2=0
+ $Y2=0
cc_130 A_N N_A_27_74#_c_158_n 0.0204399f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A_N_c_125_n N_A_27_74#_c_165_n 0.00202f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A_N_c_125_n N_A_27_74#_c_167_n 0.0119404f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_N_c_125_n N_A_27_74#_c_168_n 0.0153468f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_134 A_N N_A_27_74#_c_168_n 0.00204776f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_135 N_A_N_M1020_g N_A_27_74#_c_159_n 0.00235298f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_136 N_A_N_c_125_n N_A_27_74#_c_169_n 0.00852474f $X=0.865 $Y=1.765 $X2=0
+ $Y2=0
cc_137 A_N N_A_27_74#_c_169_n 0.0252036f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A_N_c_125_n N_A_27_74#_c_160_n 0.00550947f $X=0.865 $Y=1.765 $X2=0
+ $Y2=0
cc_139 A_N N_A_27_74#_c_160_n 0.0100197f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A_N_c_125_n N_A_27_74#_c_161_n 0.0191304f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_N_c_125_n N_A_298_368#_c_376_n 7.1556e-19 $X=0.865 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_N_c_125_n N_VPWR_c_534_n 0.0082943f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_N_c_125_n N_VPWR_c_545_n 0.00481995f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_N_c_125_n N_VPWR_c_533_n 0.00508379f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_N_M1020_g N_VGND_c_716_n 0.00495522f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_146 N_A_N_c_125_n N_VGND_c_716_n 0.0030517f $X=0.865 $Y=1.765 $X2=0 $Y2=0
cc_147 A_N N_VGND_c_716_n 0.017597f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A_N_M1020_g N_VGND_c_722_n 0.00434272f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_149 N_A_N_M1020_g N_VGND_c_731_n 0.00828717f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_150 N_A_N_M1020_g N_A_239_98#_c_808_n 0.00446029f $X=0.495 $Y=0.69 $X2=0
+ $Y2=0
cc_151 N_A_27_74#_M1018_g N_B_M1015_g 0.0160281f $X=1.985 $Y=0.81 $X2=0 $Y2=0
cc_152 N_A_27_74#_c_163_n N_B_c_245_n 0.0288123f $X=1.865 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_27_74#_c_161_n B 0.00683976f $X=1.865 $Y=1.542 $X2=0 $Y2=0
cc_154 N_A_27_74#_c_161_n N_B_c_244_n 0.0145633f $X=1.865 $Y=1.542 $X2=0 $Y2=0
cc_155 N_A_27_74#_c_162_n N_A_298_368#_c_372_n 0.00751626f $X=1.415 $Y=1.765
+ $X2=0 $Y2=0
cc_156 N_A_27_74#_c_163_n N_A_298_368#_c_372_n 0.00920205f $X=1.865 $Y=1.765
+ $X2=0 $Y2=0
cc_157 N_A_27_74#_c_163_n N_A_298_368#_c_382_n 0.0113798f $X=1.865 $Y=1.765
+ $X2=0 $Y2=0
cc_158 N_A_27_74#_c_161_n N_A_298_368#_c_382_n 0.00222461f $X=1.865 $Y=1.542
+ $X2=0 $Y2=0
cc_159 N_A_27_74#_c_163_n N_A_298_368#_c_373_n 6.39089e-19 $X=1.865 $Y=1.765
+ $X2=0 $Y2=0
cc_160 N_A_27_74#_c_162_n N_A_298_368#_c_376_n 0.00501186f $X=1.415 $Y=1.765
+ $X2=0 $Y2=0
cc_161 N_A_27_74#_c_163_n N_A_298_368#_c_376_n 0.00813193f $X=1.865 $Y=1.765
+ $X2=0 $Y2=0
cc_162 N_A_27_74#_c_167_n N_A_298_368#_c_376_n 0.00409238f $X=0.64 $Y=1.985
+ $X2=0 $Y2=0
cc_163 N_A_27_74#_c_160_n N_A_298_368#_c_376_n 0.00613533f $X=1.36 $Y=1.485
+ $X2=0 $Y2=0
cc_164 N_A_27_74#_c_161_n N_A_298_368#_c_376_n 0.00872242f $X=1.865 $Y=1.542
+ $X2=0 $Y2=0
cc_165 N_A_27_74#_c_162_n N_A_298_368#_c_362_n 4.11163e-19 $X=1.415 $Y=1.765
+ $X2=0 $Y2=0
cc_166 N_A_27_74#_M1000_g N_A_298_368#_c_362_n 0.00398237f $X=1.555 $Y=0.81
+ $X2=0 $Y2=0
cc_167 N_A_27_74#_c_163_n N_A_298_368#_c_362_n 0.00142212f $X=1.865 $Y=1.765
+ $X2=0 $Y2=0
cc_168 N_A_27_74#_c_160_n N_A_298_368#_c_362_n 0.0318758f $X=1.36 $Y=1.485 $X2=0
+ $Y2=0
cc_169 N_A_27_74#_c_161_n N_A_298_368#_c_362_n 0.0212189f $X=1.865 $Y=1.542
+ $X2=0 $Y2=0
cc_170 N_A_27_74#_M1000_g N_A_298_368#_c_363_n 7.50786e-19 $X=1.555 $Y=0.81
+ $X2=0 $Y2=0
cc_171 N_A_27_74#_M1018_g N_A_298_368#_c_363_n 0.00453293f $X=1.985 $Y=0.81
+ $X2=0 $Y2=0
cc_172 N_A_27_74#_c_168_n N_VPWR_M1010_d 0.00145634f $X=1.135 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_27_74#_c_160_n N_VPWR_M1010_d 0.00170732f $X=1.36 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_27_74#_c_162_n N_VPWR_c_534_n 0.00689359f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A_27_74#_c_167_n N_VPWR_c_534_n 0.0323093f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_27_74#_c_168_n N_VPWR_c_534_n 0.011191f $X=1.135 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_27_74#_c_160_n N_VPWR_c_534_n 0.0131018f $X=1.36 $Y=1.485 $X2=0 $Y2=0
cc_178 N_A_27_74#_c_161_n N_VPWR_c_534_n 5.00418e-19 $X=1.865 $Y=1.542 $X2=0
+ $Y2=0
cc_179 N_A_27_74#_c_163_n N_VPWR_c_535_n 0.00528632f $X=1.865 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A_27_74#_c_167_n N_VPWR_c_545_n 0.0097982f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_27_74#_c_162_n N_VPWR_c_546_n 0.00481995f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_27_74#_c_163_n N_VPWR_c_546_n 0.00481995f $X=1.865 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_27_74#_c_162_n N_VPWR_c_533_n 0.00508379f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A_27_74#_c_163_n N_VPWR_c_533_n 0.00508379f $X=1.865 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_27_74#_c_167_n N_VPWR_c_533_n 0.0111907f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_27_74#_M1000_g N_VGND_c_716_n 0.00147712f $X=1.555 $Y=0.81 $X2=0
+ $Y2=0
cc_187 N_A_27_74#_c_157_n N_VGND_c_716_n 0.0254897f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_188 N_A_27_74#_c_168_n N_VGND_c_716_n 0.00107831f $X=1.135 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A_27_74#_c_157_n N_VGND_c_722_n 0.0145488f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_190 N_A_27_74#_M1000_g N_VGND_c_723_n 7.4413e-19 $X=1.555 $Y=0.81 $X2=0 $Y2=0
cc_191 N_A_27_74#_M1018_g N_VGND_c_723_n 7.21231e-19 $X=1.985 $Y=0.81 $X2=0
+ $Y2=0
cc_192 N_A_27_74#_c_157_n N_VGND_c_731_n 0.0119924f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_193 N_A_27_74#_M1000_g N_A_239_98#_c_808_n 0.0106946f $X=1.555 $Y=0.81 $X2=0
+ $Y2=0
cc_194 N_A_27_74#_M1018_g N_A_239_98#_c_808_n 6.65289e-19 $X=1.985 $Y=0.81 $X2=0
+ $Y2=0
cc_195 N_A_27_74#_c_160_n N_A_239_98#_c_808_n 0.0281374f $X=1.36 $Y=1.485 $X2=0
+ $Y2=0
cc_196 N_A_27_74#_c_161_n N_A_239_98#_c_808_n 0.00224193f $X=1.865 $Y=1.542
+ $X2=0 $Y2=0
cc_197 N_A_27_74#_M1000_g N_A_239_98#_c_809_n 0.00902186f $X=1.555 $Y=0.81 $X2=0
+ $Y2=0
cc_198 N_A_27_74#_M1018_g N_A_239_98#_c_809_n 0.00927815f $X=1.985 $Y=0.81 $X2=0
+ $Y2=0
cc_199 N_A_27_74#_M1000_g N_A_239_98#_c_810_n 0.00187523f $X=1.555 $Y=0.81 $X2=0
+ $Y2=0
cc_200 N_A_27_74#_M1000_g N_A_239_98#_c_812_n 6.91231e-19 $X=1.555 $Y=0.81 $X2=0
+ $Y2=0
cc_201 N_A_27_74#_M1018_g N_A_239_98#_c_812_n 0.00647313f $X=1.985 $Y=0.81 $X2=0
+ $Y2=0
cc_202 N_A_27_74#_M1018_g N_A_239_98#_c_813_n 0.00521983f $X=1.985 $Y=0.81 $X2=0
+ $Y2=0
cc_203 N_B_c_246_n N_C_c_302_n 0.0246387f $X=2.865 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_204 N_B_M1016_g N_C_c_299_n 0.0178135f $X=2.915 $Y=0.81 $X2=0 $Y2=0
cc_205 B N_C_c_299_n 2.20256e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_206 N_B_c_244_n N_C_c_299_n 0.0100708f $X=2.865 $Y=1.557 $X2=0 $Y2=0
cc_207 B N_C_c_301_n 0.0286185f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_208 N_B_c_244_n N_C_c_301_n 0.00463881f $X=2.865 $Y=1.557 $X2=0 $Y2=0
cc_209 N_B_c_245_n N_A_298_368#_c_372_n 6.39089e-19 $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_210 N_B_c_245_n N_A_298_368#_c_382_n 0.0124513f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_211 B N_A_298_368#_c_382_n 0.0312432f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_212 N_B_c_245_n N_A_298_368#_c_373_n 0.00920205f $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_B_c_246_n N_A_298_368#_c_373_n 0.00935377f $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_B_c_246_n N_A_298_368#_c_402_n 0.0167844f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_215 N_B_c_246_n N_A_298_368#_c_374_n 8.78039e-19 $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_216 N_B_c_245_n N_A_298_368#_c_362_n 8.71714e-19 $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_217 B N_A_298_368#_c_362_n 0.0326263f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_218 N_B_c_244_n N_A_298_368#_c_362_n 2.96541e-19 $X=2.865 $Y=1.557 $X2=0
+ $Y2=0
cc_219 N_B_c_245_n N_A_298_368#_c_407_n 4.27055e-19 $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_220 N_B_c_246_n N_A_298_368#_c_407_n 9.50925e-19 $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_221 B N_A_298_368#_c_407_n 0.0210582f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_222 N_B_c_244_n N_A_298_368#_c_407_n 0.00137486f $X=2.865 $Y=1.557 $X2=0
+ $Y2=0
cc_223 N_B_c_245_n N_VPWR_c_535_n 0.00528632f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_224 N_B_c_246_n N_VPWR_c_536_n 0.00577667f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_225 N_B_c_245_n N_VPWR_c_547_n 0.00481995f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_226 N_B_c_246_n N_VPWR_c_547_n 0.00481995f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_227 N_B_c_245_n N_VPWR_c_533_n 0.00508379f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_228 N_B_c_246_n N_VPWR_c_533_n 0.00508379f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_229 N_B_M1016_g N_VGND_c_717_n 0.00506675f $X=2.915 $Y=0.81 $X2=0 $Y2=0
cc_230 N_B_M1015_g N_VGND_c_723_n 0.00319047f $X=2.415 $Y=0.81 $X2=0 $Y2=0
cc_231 N_B_M1016_g N_VGND_c_723_n 0.00364981f $X=2.915 $Y=0.81 $X2=0 $Y2=0
cc_232 N_B_M1015_g N_VGND_c_731_n 0.00427039f $X=2.415 $Y=0.81 $X2=0 $Y2=0
cc_233 N_B_M1016_g N_VGND_c_731_n 0.00508379f $X=2.915 $Y=0.81 $X2=0 $Y2=0
cc_234 N_B_M1015_g N_A_239_98#_c_811_n 0.0123579f $X=2.415 $Y=0.81 $X2=0 $Y2=0
cc_235 N_B_M1016_g N_A_239_98#_c_811_n 0.0119434f $X=2.915 $Y=0.81 $X2=0 $Y2=0
cc_236 B N_A_239_98#_c_811_n 0.00376415f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_237 N_B_M1015_g N_A_239_98#_c_812_n 0.00534802f $X=2.415 $Y=0.81 $X2=0 $Y2=0
cc_238 N_B_M1016_g N_A_239_98#_c_812_n 0.00119972f $X=2.915 $Y=0.81 $X2=0 $Y2=0
cc_239 N_B_M1015_g N_A_239_98#_c_813_n 0.00652109f $X=2.415 $Y=0.81 $X2=0 $Y2=0
cc_240 B N_A_239_98#_c_813_n 0.0252291f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B_c_244_n N_A_239_98#_c_813_n 3.5991e-19 $X=2.865 $Y=1.557 $X2=0 $Y2=0
cc_242 N_B_M1016_g N_A_498_98#_c_853_n 0.014257f $X=2.915 $Y=0.81 $X2=0 $Y2=0
cc_243 N_B_M1015_g N_A_498_98#_c_855_n 0.00188875f $X=2.415 $Y=0.81 $X2=0 $Y2=0
cc_244 N_B_M1016_g N_A_498_98#_c_855_n 0.00818413f $X=2.915 $Y=0.81 $X2=0 $Y2=0
cc_245 B N_A_498_98#_c_855_n 0.0175828f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_246 N_B_c_244_n N_A_498_98#_c_855_n 0.00386322f $X=2.865 $Y=1.557 $X2=0 $Y2=0
cc_247 N_C_c_303_n N_A_298_368#_c_366_n 0.022126f $X=3.925 $Y=1.765 $X2=0 $Y2=0
cc_248 N_C_c_299_n N_A_298_368#_c_356_n 0.00588736f $X=4.015 $Y=1.28 $X2=0 $Y2=0
cc_249 N_C_c_300_n N_A_298_368#_M1006_g 0.0183935f $X=4.335 $Y=1.205 $X2=0 $Y2=0
cc_250 N_C_c_302_n N_A_298_368#_c_373_n 8.46192e-19 $X=3.475 $Y=1.765 $X2=0
+ $Y2=0
cc_251 N_C_c_302_n N_A_298_368#_c_402_n 0.0126919f $X=3.475 $Y=1.765 $X2=0 $Y2=0
cc_252 N_C_c_299_n N_A_298_368#_c_402_n 7.64221e-19 $X=4.015 $Y=1.28 $X2=0 $Y2=0
cc_253 N_C_c_301_n N_A_298_368#_c_402_n 0.0392083f $X=3.395 $Y=1.515 $X2=0 $Y2=0
cc_254 N_C_c_302_n N_A_298_368#_c_374_n 0.0102214f $X=3.475 $Y=1.765 $X2=0 $Y2=0
cc_255 N_C_c_303_n N_A_298_368#_c_374_n 0.00975269f $X=3.925 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_C_c_302_n N_A_298_368#_c_375_n 0.00317149f $X=3.475 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_C_c_303_n N_A_298_368#_c_375_n 0.00323388f $X=3.925 $Y=1.765 $X2=0
+ $Y2=0
cc_258 N_C_c_299_n N_A_298_368#_c_375_n 0.00810591f $X=4.015 $Y=1.28 $X2=0 $Y2=0
cc_259 N_C_c_301_n N_A_298_368#_c_375_n 0.0115569f $X=3.395 $Y=1.515 $X2=0 $Y2=0
cc_260 N_C_c_299_n N_A_298_368#_c_424_n 0.00792271f $X=4.015 $Y=1.28 $X2=0 $Y2=0
cc_261 N_C_c_301_n N_A_298_368#_c_424_n 0.0141716f $X=3.395 $Y=1.515 $X2=0 $Y2=0
cc_262 N_C_c_298_n N_A_298_368#_c_361_n 3.87319e-19 $X=4.26 $Y=1.28 $X2=0 $Y2=0
cc_263 N_C_c_302_n N_A_298_368#_c_427_n 4.27055e-19 $X=3.475 $Y=1.765 $X2=0
+ $Y2=0
cc_264 N_C_c_303_n N_A_298_368#_c_427_n 0.00205145f $X=3.925 $Y=1.765 $X2=0
+ $Y2=0
cc_265 N_C_c_299_n N_A_298_368#_c_427_n 0.00593494f $X=4.015 $Y=1.28 $X2=0 $Y2=0
cc_266 N_C_c_301_n N_A_298_368#_c_427_n 0.00161377f $X=3.395 $Y=1.515 $X2=0
+ $Y2=0
cc_267 N_C_c_298_n N_A_298_368#_c_364_n 0.0127946f $X=4.26 $Y=1.28 $X2=0 $Y2=0
cc_268 N_C_c_299_n N_A_298_368#_c_364_n 0.0127038f $X=4.015 $Y=1.28 $X2=0 $Y2=0
cc_269 N_C_c_298_n N_A_298_368#_c_365_n 0.00199908f $X=4.26 $Y=1.28 $X2=0 $Y2=0
cc_270 N_C_c_302_n N_VPWR_c_536_n 0.00867226f $X=3.475 $Y=1.765 $X2=0 $Y2=0
cc_271 N_C_c_302_n N_VPWR_c_537_n 0.00481995f $X=3.475 $Y=1.765 $X2=0 $Y2=0
cc_272 N_C_c_303_n N_VPWR_c_537_n 0.00451858f $X=3.925 $Y=1.765 $X2=0 $Y2=0
cc_273 N_C_c_303_n N_VPWR_c_538_n 0.0125738f $X=3.925 $Y=1.765 $X2=0 $Y2=0
cc_274 N_C_c_302_n N_VPWR_c_533_n 0.00508379f $X=3.475 $Y=1.765 $X2=0 $Y2=0
cc_275 N_C_c_303_n N_VPWR_c_533_n 0.00508379f $X=3.925 $Y=1.765 $X2=0 $Y2=0
cc_276 N_C_c_297_n N_VGND_c_717_n 0.00974237f $X=3.905 $Y=1.205 $X2=0 $Y2=0
cc_277 N_C_c_300_n N_VGND_c_717_n 4.59889e-19 $X=4.335 $Y=1.205 $X2=0 $Y2=0
cc_278 N_C_c_300_n N_VGND_c_718_n 0.00531636f $X=4.335 $Y=1.205 $X2=0 $Y2=0
cc_279 N_C_c_297_n N_VGND_c_724_n 0.00421418f $X=3.905 $Y=1.205 $X2=0 $Y2=0
cc_280 N_C_c_300_n N_VGND_c_724_n 0.00485498f $X=4.335 $Y=1.205 $X2=0 $Y2=0
cc_281 N_C_c_297_n N_VGND_c_731_n 0.00432128f $X=3.905 $Y=1.205 $X2=0 $Y2=0
cc_282 N_C_c_300_n N_VGND_c_731_n 0.00514438f $X=4.335 $Y=1.205 $X2=0 $Y2=0
cc_283 N_C_c_297_n N_A_239_98#_c_811_n 5.33566e-19 $X=3.905 $Y=1.205 $X2=0 $Y2=0
cc_284 N_C_c_297_n N_A_498_98#_c_853_n 0.0155958f $X=3.905 $Y=1.205 $X2=0 $Y2=0
cc_285 N_C_c_298_n N_A_498_98#_c_853_n 0.00262633f $X=4.26 $Y=1.28 $X2=0 $Y2=0
cc_286 N_C_c_299_n N_A_498_98#_c_853_n 0.0207597f $X=4.015 $Y=1.28 $X2=0 $Y2=0
cc_287 N_C_c_300_n N_A_498_98#_c_853_n 0.00345767f $X=4.335 $Y=1.205 $X2=0 $Y2=0
cc_288 N_C_c_301_n N_A_498_98#_c_853_n 0.0435313f $X=3.395 $Y=1.515 $X2=0 $Y2=0
cc_289 N_C_c_300_n N_A_498_98#_c_854_n 0.00632016f $X=4.335 $Y=1.205 $X2=0 $Y2=0
cc_290 N_A_298_368#_c_382_n N_VPWR_M1008_s 0.00665611f $X=2.475 $Y=2.035 $X2=0
+ $Y2=0
cc_291 N_A_298_368#_c_402_n N_VPWR_M1007_s 0.00936632f $X=3.535 $Y=2.035 $X2=0
+ $Y2=0
cc_292 N_A_298_368#_c_376_n N_VPWR_c_534_n 0.0323689f $X=1.64 $Y=1.985 $X2=0
+ $Y2=0
cc_293 N_A_298_368#_c_372_n N_VPWR_c_535_n 0.0221782f $X=1.64 $Y=2.695 $X2=0
+ $Y2=0
cc_294 N_A_298_368#_c_382_n N_VPWR_c_535_n 0.0232685f $X=2.475 $Y=2.035 $X2=0
+ $Y2=0
cc_295 N_A_298_368#_c_373_n N_VPWR_c_535_n 0.0221782f $X=2.64 $Y=2.715 $X2=0
+ $Y2=0
cc_296 N_A_298_368#_c_373_n N_VPWR_c_536_n 0.0221782f $X=2.64 $Y=2.715 $X2=0
+ $Y2=0
cc_297 N_A_298_368#_c_402_n N_VPWR_c_536_n 0.0249771f $X=3.535 $Y=2.035 $X2=0
+ $Y2=0
cc_298 N_A_298_368#_c_374_n N_VPWR_c_536_n 0.0353739f $X=3.7 $Y=2.715 $X2=0
+ $Y2=0
cc_299 N_A_298_368#_c_374_n N_VPWR_c_537_n 0.0107215f $X=3.7 $Y=2.715 $X2=0
+ $Y2=0
cc_300 N_A_298_368#_c_366_n N_VPWR_c_538_n 0.010964f $X=4.51 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_298_368#_c_374_n N_VPWR_c_538_n 0.0578659f $X=3.7 $Y=2.715 $X2=0
+ $Y2=0
cc_302 N_A_298_368#_c_375_n N_VPWR_c_538_n 0.00961521f $X=3.815 $Y=1.95 $X2=0
+ $Y2=0
cc_303 N_A_298_368#_c_427_n N_VPWR_c_538_n 0.0140085f $X=3.7 $Y=2.035 $X2=0
+ $Y2=0
cc_304 N_A_298_368#_c_364_n N_VPWR_c_538_n 0.0256059f $X=4.755 $Y=1.465 $X2=0
+ $Y2=0
cc_305 N_A_298_368#_c_369_n N_VPWR_c_539_n 0.00687925f $X=4.96 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_298_368#_c_370_n N_VPWR_c_539_n 0.00687925f $X=5.51 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_298_368#_c_371_n N_VPWR_c_540_n 0.0198182f $X=5.96 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_A_298_368#_c_365_n N_VPWR_c_540_n 3.20042e-19 $X=5.96 $Y=1.532 $X2=0
+ $Y2=0
cc_309 N_A_298_368#_c_366_n N_VPWR_c_541_n 0.00445602f $X=4.51 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_A_298_368#_c_369_n N_VPWR_c_541_n 0.00445602f $X=4.96 $Y=1.765 $X2=0
+ $Y2=0
cc_311 N_A_298_368#_c_370_n N_VPWR_c_543_n 0.00445602f $X=5.51 $Y=1.765 $X2=0
+ $Y2=0
cc_312 N_A_298_368#_c_371_n N_VPWR_c_543_n 0.00445602f $X=5.96 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_A_298_368#_c_372_n N_VPWR_c_546_n 0.00976219f $X=1.64 $Y=2.695 $X2=0
+ $Y2=0
cc_314 N_A_298_368#_c_373_n N_VPWR_c_547_n 0.00976219f $X=2.64 $Y=2.715 $X2=0
+ $Y2=0
cc_315 N_A_298_368#_c_366_n N_VPWR_c_533_n 0.00861719f $X=4.51 $Y=1.765 $X2=0
+ $Y2=0
cc_316 N_A_298_368#_c_369_n N_VPWR_c_533_n 0.00857797f $X=4.96 $Y=1.765 $X2=0
+ $Y2=0
cc_317 N_A_298_368#_c_370_n N_VPWR_c_533_n 0.00857797f $X=5.51 $Y=1.765 $X2=0
+ $Y2=0
cc_318 N_A_298_368#_c_371_n N_VPWR_c_533_n 0.00861002f $X=5.96 $Y=1.765 $X2=0
+ $Y2=0
cc_319 N_A_298_368#_c_372_n N_VPWR_c_533_n 0.0111764f $X=1.64 $Y=2.695 $X2=0
+ $Y2=0
cc_320 N_A_298_368#_c_373_n N_VPWR_c_533_n 0.0111764f $X=2.64 $Y=2.715 $X2=0
+ $Y2=0
cc_321 N_A_298_368#_c_374_n N_VPWR_c_533_n 0.0123362f $X=3.7 $Y=2.715 $X2=0
+ $Y2=0
cc_322 N_A_298_368#_c_366_n N_X_c_638_n 0.0107529f $X=4.51 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A_298_368#_c_369_n N_X_c_638_n 0.0123916f $X=4.96 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A_298_368#_c_370_n N_X_c_638_n 6.94077e-19 $X=5.51 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A_298_368#_c_369_n N_X_c_639_n 0.0125195f $X=4.96 $Y=1.765 $X2=0 $Y2=0
cc_326 N_A_298_368#_c_370_n N_X_c_639_n 0.0125195f $X=5.51 $Y=1.765 $X2=0 $Y2=0
cc_327 N_A_298_368#_c_361_n N_X_c_639_n 0.0492346f $X=4.92 $Y=1.465 $X2=0 $Y2=0
cc_328 N_A_298_368#_c_365_n N_X_c_639_n 0.0116817f $X=5.96 $Y=1.532 $X2=0 $Y2=0
cc_329 N_A_298_368#_c_366_n N_X_c_640_n 0.00256459f $X=4.51 $Y=1.765 $X2=0 $Y2=0
cc_330 N_A_298_368#_c_355_n N_X_c_640_n 0.00708737f $X=4.755 $Y=1.67 $X2=0 $Y2=0
cc_331 N_A_298_368#_c_356_n N_X_c_640_n 3.62994e-19 $X=4.6 $Y=1.67 $X2=0 $Y2=0
cc_332 N_A_298_368#_c_369_n N_X_c_640_n 9.3899e-19 $X=4.96 $Y=1.765 $X2=0 $Y2=0
cc_333 N_A_298_368#_c_375_n N_X_c_640_n 4.82305e-19 $X=3.815 $Y=1.95 $X2=0 $Y2=0
cc_334 N_A_298_368#_c_364_n N_X_c_640_n 0.0269477f $X=4.755 $Y=1.465 $X2=0 $Y2=0
cc_335 N_A_298_368#_c_365_n N_X_c_640_n 4.80986e-19 $X=5.96 $Y=1.532 $X2=0 $Y2=0
cc_336 N_A_298_368#_M1006_g N_X_c_631_n 0.00323888f $X=4.845 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A_298_368#_M1011_g N_X_c_631_n 4.69391e-19 $X=5.345 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A_298_368#_M1011_g N_X_c_632_n 0.0125602f $X=5.345 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A_298_368#_M1013_g N_X_c_632_n 0.0144374f $X=5.795 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A_298_368#_c_484_p N_X_c_632_n 0.0405722f $X=5.6 $Y=1.465 $X2=0 $Y2=0
cc_341 N_A_298_368#_c_365_n N_X_c_632_n 0.00305348f $X=5.96 $Y=1.532 $X2=0 $Y2=0
cc_342 N_A_298_368#_M1006_g N_X_c_633_n 9.62947e-19 $X=4.845 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A_298_368#_c_484_p N_X_c_633_n 0.0210849f $X=5.6 $Y=1.465 $X2=0 $Y2=0
cc_344 N_A_298_368#_c_365_n N_X_c_633_n 0.00426938f $X=5.96 $Y=1.532 $X2=0 $Y2=0
cc_345 N_A_298_368#_c_369_n N_X_c_641_n 6.94077e-19 $X=4.96 $Y=1.765 $X2=0 $Y2=0
cc_346 N_A_298_368#_c_370_n N_X_c_641_n 0.0123916f $X=5.51 $Y=1.765 $X2=0 $Y2=0
cc_347 N_A_298_368#_c_371_n N_X_c_641_n 0.0165744f $X=5.96 $Y=1.765 $X2=0 $Y2=0
cc_348 N_A_298_368#_M1013_g N_X_c_634_n 3.98709e-19 $X=5.795 $Y=0.74 $X2=0 $Y2=0
cc_349 N_A_298_368#_M1017_g N_X_c_634_n 3.98398e-19 $X=6.225 $Y=0.74 $X2=0 $Y2=0
cc_350 N_A_298_368#_M1013_g N_X_c_635_n 0.00398237f $X=5.795 $Y=0.74 $X2=0 $Y2=0
cc_351 N_A_298_368#_c_371_n N_X_c_635_n 0.00127528f $X=5.96 $Y=1.765 $X2=0 $Y2=0
cc_352 N_A_298_368#_M1017_g N_X_c_635_n 0.00408495f $X=6.225 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A_298_368#_c_484_p N_X_c_635_n 0.0249855f $X=5.6 $Y=1.465 $X2=0 $Y2=0
cc_354 N_A_298_368#_c_365_n N_X_c_635_n 0.0303553f $X=5.96 $Y=1.532 $X2=0 $Y2=0
cc_355 N_A_298_368#_c_365_n N_X_c_643_n 0.00644978f $X=5.96 $Y=1.532 $X2=0 $Y2=0
cc_356 N_A_298_368#_c_370_n N_X_c_644_n 9.3899e-19 $X=5.51 $Y=1.765 $X2=0 $Y2=0
cc_357 N_A_298_368#_c_371_n N_X_c_644_n 0.0144489f $X=5.96 $Y=1.765 $X2=0 $Y2=0
cc_358 N_A_298_368#_c_484_p N_X_c_644_n 0.0163751f $X=5.6 $Y=1.465 $X2=0 $Y2=0
cc_359 N_A_298_368#_c_365_n N_X_c_644_n 0.0103015f $X=5.96 $Y=1.532 $X2=0 $Y2=0
cc_360 N_A_298_368#_c_371_n X 7.93392e-19 $X=5.96 $Y=1.765 $X2=0 $Y2=0
cc_361 N_A_298_368#_c_365_n X 0.00125888f $X=5.96 $Y=1.532 $X2=0 $Y2=0
cc_362 N_A_298_368#_c_356_n N_VGND_c_718_n 0.00163829f $X=4.6 $Y=1.67 $X2=0
+ $Y2=0
cc_363 N_A_298_368#_M1006_g N_VGND_c_718_n 0.0142051f $X=4.845 $Y=0.74 $X2=0
+ $Y2=0
cc_364 N_A_298_368#_M1011_g N_VGND_c_718_n 5.30714e-19 $X=5.345 $Y=0.74 $X2=0
+ $Y2=0
cc_365 N_A_298_368#_c_361_n N_VGND_c_718_n 0.00318079f $X=4.92 $Y=1.465 $X2=0
+ $Y2=0
cc_366 N_A_298_368#_c_364_n N_VGND_c_718_n 0.0153656f $X=4.755 $Y=1.465 $X2=0
+ $Y2=0
cc_367 N_A_298_368#_c_365_n N_VGND_c_718_n 3.70873e-19 $X=5.96 $Y=1.532 $X2=0
+ $Y2=0
cc_368 N_A_298_368#_M1006_g N_VGND_c_719_n 4.47887e-19 $X=4.845 $Y=0.74 $X2=0
+ $Y2=0
cc_369 N_A_298_368#_M1011_g N_VGND_c_719_n 0.009906f $X=5.345 $Y=0.74 $X2=0
+ $Y2=0
cc_370 N_A_298_368#_M1013_g N_VGND_c_719_n 0.00834923f $X=5.795 $Y=0.74 $X2=0
+ $Y2=0
cc_371 N_A_298_368#_M1017_g N_VGND_c_719_n 4.52684e-19 $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_372 N_A_298_368#_M1013_g N_VGND_c_721_n 5.57023e-19 $X=5.795 $Y=0.74 $X2=0
+ $Y2=0
cc_373 N_A_298_368#_M1017_g N_VGND_c_721_n 0.0150765f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_374 N_A_298_368#_M1006_g N_VGND_c_725_n 0.00383152f $X=4.845 $Y=0.74 $X2=0
+ $Y2=0
cc_375 N_A_298_368#_M1011_g N_VGND_c_725_n 0.00383152f $X=5.345 $Y=0.74 $X2=0
+ $Y2=0
cc_376 N_A_298_368#_M1013_g N_VGND_c_726_n 0.00444681f $X=5.795 $Y=0.74 $X2=0
+ $Y2=0
cc_377 N_A_298_368#_M1017_g N_VGND_c_726_n 0.00383152f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_378 N_A_298_368#_M1006_g N_VGND_c_731_n 0.00758198f $X=4.845 $Y=0.74 $X2=0
+ $Y2=0
cc_379 N_A_298_368#_M1011_g N_VGND_c_731_n 0.00758198f $X=5.345 $Y=0.74 $X2=0
+ $Y2=0
cc_380 N_A_298_368#_M1013_g N_VGND_c_731_n 0.00877518f $X=5.795 $Y=0.74 $X2=0
+ $Y2=0
cc_381 N_A_298_368#_M1017_g N_VGND_c_731_n 0.0075754f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_382 N_A_298_368#_c_363_n N_A_239_98#_c_808_n 0.0205845f $X=1.775 $Y=1.15
+ $X2=0 $Y2=0
cc_383 N_A_298_368#_c_527_p N_A_239_98#_c_809_n 0.0133f $X=1.77 $Y=0.87 $X2=0
+ $Y2=0
cc_384 N_A_298_368#_c_363_n N_A_239_98#_c_812_n 0.0215085f $X=1.775 $Y=1.15
+ $X2=0 $Y2=0
cc_385 N_A_298_368#_M1006_g N_A_498_98#_c_853_n 2.71064e-19 $X=4.845 $Y=0.74
+ $X2=0 $Y2=0
cc_386 N_A_298_368#_c_424_n N_A_498_98#_c_853_n 0.00905654f $X=3.9 $Y=1.545
+ $X2=0 $Y2=0
cc_387 N_A_298_368#_c_364_n N_A_498_98#_c_853_n 0.0211484f $X=4.755 $Y=1.465
+ $X2=0 $Y2=0
cc_388 N_A_298_368#_c_362_n N_A_498_98#_c_855_n 8.78562e-19 $X=1.67 $Y=1.82
+ $X2=0 $Y2=0
cc_389 N_VPWR_c_538_n N_X_c_638_n 0.0386506f $X=4.235 $Y=1.985 $X2=0 $Y2=0
cc_390 N_VPWR_c_539_n N_X_c_638_n 0.0323093f $X=5.235 $Y=2.25 $X2=0 $Y2=0
cc_391 N_VPWR_c_541_n N_X_c_638_n 0.014552f $X=5.07 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_c_533_n N_X_c_638_n 0.0119791f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_393 N_VPWR_M1005_s N_X_c_639_n 0.00332584f $X=5.035 $Y=1.84 $X2=0 $Y2=0
cc_394 N_VPWR_c_539_n N_X_c_639_n 0.0232685f $X=5.235 $Y=2.25 $X2=0 $Y2=0
cc_395 N_VPWR_c_538_n N_X_c_640_n 0.00711242f $X=4.235 $Y=1.985 $X2=0 $Y2=0
cc_396 N_VPWR_c_539_n N_X_c_641_n 0.0323093f $X=5.235 $Y=2.25 $X2=0 $Y2=0
cc_397 N_VPWR_c_540_n N_X_c_641_n 0.0323093f $X=6.235 $Y=2.25 $X2=0 $Y2=0
cc_398 N_VPWR_c_543_n N_X_c_641_n 0.014552f $X=6.07 $Y=3.33 $X2=0 $Y2=0
cc_399 N_VPWR_c_533_n N_X_c_641_n 0.0119791f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_400 N_VPWR_M1012_s N_X_c_643_n 0.00411851f $X=6.035 $Y=1.84 $X2=0 $Y2=0
cc_401 N_VPWR_c_540_n N_X_c_643_n 0.0211167f $X=6.235 $Y=2.25 $X2=0 $Y2=0
cc_402 N_VPWR_c_540_n N_X_c_644_n 0.0011721f $X=6.235 $Y=2.25 $X2=0 $Y2=0
cc_403 N_VPWR_M1012_s X 5.82949e-19 $X=6.035 $Y=1.84 $X2=0 $Y2=0
cc_404 N_VPWR_c_540_n X 0.00293678f $X=6.235 $Y=2.25 $X2=0 $Y2=0
cc_405 N_X_c_632_n N_VGND_M1011_d 0.00197722f $X=5.925 $Y=1.045 $X2=0 $Y2=0
cc_406 N_X_c_631_n N_VGND_c_718_n 0.0236466f $X=5.13 $Y=0.515 $X2=0 $Y2=0
cc_407 N_X_c_633_n N_VGND_c_718_n 0.00729487f $X=5.215 $Y=1.045 $X2=0 $Y2=0
cc_408 N_X_c_631_n N_VGND_c_719_n 0.0164981f $X=5.13 $Y=0.515 $X2=0 $Y2=0
cc_409 N_X_c_632_n N_VGND_c_719_n 0.0171813f $X=5.925 $Y=1.045 $X2=0 $Y2=0
cc_410 N_X_c_634_n N_VGND_c_719_n 0.0151391f $X=6.01 $Y=0.515 $X2=0 $Y2=0
cc_411 N_X_c_634_n N_VGND_c_721_n 0.0236097f $X=6.01 $Y=0.515 $X2=0 $Y2=0
cc_412 N_X_c_643_n N_VGND_c_721_n 0.0027645f $X=6.365 $Y=1.885 $X2=0 $Y2=0
cc_413 N_X_c_636_n N_VGND_c_721_n 0.00729487f $X=6.015 $Y=1.045 $X2=0 $Y2=0
cc_414 X N_VGND_c_721_n 0.0109822f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_415 N_X_c_631_n N_VGND_c_725_n 0.011066f $X=5.13 $Y=0.515 $X2=0 $Y2=0
cc_416 N_X_c_634_n N_VGND_c_726_n 0.00794252f $X=6.01 $Y=0.515 $X2=0 $Y2=0
cc_417 N_X_c_631_n N_VGND_c_731_n 0.00915947f $X=5.13 $Y=0.515 $X2=0 $Y2=0
cc_418 N_X_c_634_n N_VGND_c_731_n 0.00657413f $X=6.01 $Y=0.515 $X2=0 $Y2=0
cc_419 N_VGND_c_716_n N_A_239_98#_c_808_n 0.0322448f $X=0.71 $Y=0.495 $X2=0
+ $Y2=0
cc_420 N_VGND_c_723_n N_A_239_98#_c_809_n 0.0341126f $X=3.525 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_731_n N_A_239_98#_c_809_n 0.0199228f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_716_n N_A_239_98#_c_810_n 0.00995436f $X=0.71 $Y=0.495 $X2=0
+ $Y2=0
cc_423 N_VGND_c_723_n N_A_239_98#_c_810_n 0.0236566f $X=3.525 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_731_n N_A_239_98#_c_810_n 0.0128296f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_717_n N_A_239_98#_c_811_n 0.0177417f $X=3.69 $Y=0.675 $X2=0
+ $Y2=0
cc_426 N_VGND_c_723_n N_A_239_98#_c_811_n 0.0253003f $X=3.525 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_731_n N_A_239_98#_c_811_n 0.0302919f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_c_723_n N_A_239_98#_c_812_n 0.0235133f $X=3.525 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_731_n N_A_239_98#_c_812_n 0.0127519f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_M1003_s N_A_498_98#_c_853_n 0.00299905f $X=3.545 $Y=0.47 $X2=0
+ $Y2=0
cc_431 N_VGND_c_717_n N_A_498_98#_c_853_n 0.0219405f $X=3.69 $Y=0.675 $X2=0
+ $Y2=0
cc_432 N_VGND_c_718_n N_A_498_98#_c_853_n 0.00558932f $X=4.63 $Y=0.515 $X2=0
+ $Y2=0
cc_433 N_VGND_c_717_n N_A_498_98#_c_854_n 0.0147061f $X=3.69 $Y=0.675 $X2=0
+ $Y2=0
cc_434 N_VGND_c_718_n N_A_498_98#_c_854_n 0.01996f $X=4.63 $Y=0.515 $X2=0 $Y2=0
cc_435 N_VGND_c_724_n N_A_498_98#_c_854_n 0.0078096f $X=4.465 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_731_n N_A_498_98#_c_854_n 0.0085649f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_437 N_A_239_98#_c_811_n N_A_498_98#_M1015_s 0.00239464f $X=3.13 $Y=0.635
+ $X2=-0.19 $Y2=-0.245
cc_438 N_A_239_98#_M1016_d N_A_498_98#_c_853_n 0.0037934f $X=2.99 $Y=0.49 $X2=0
+ $Y2=0
cc_439 N_A_239_98#_c_811_n N_A_498_98#_c_853_n 0.0182583f $X=3.13 $Y=0.635 $X2=0
+ $Y2=0
cc_440 N_A_239_98#_c_811_n N_A_498_98#_c_855_n 0.020173f $X=3.13 $Y=0.635 $X2=0
+ $Y2=0
cc_441 N_A_239_98#_c_813_n N_A_498_98#_c_855_n 0.0105463f $X=2.2 $Y=0.635 $X2=0
+ $Y2=0
