* File: sky130_fd_sc_hs__or3_2.spice
* Created: Thu Aug 27 21:05:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__or3_2.pex.spice"
.subckt sky130_fd_sc_hs__or3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_C_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1616 AS=0.1824 PD=1.145 PS=1.85 NRD=20.616 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_27_74#_M1008_d N_B_M1008_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.1616 PD=0.99 PS=1.145 NRD=0 NRS=21.552 M=1 R=4.26667 SA=75000.9
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_27_74#_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.179293 AS=0.112 PD=1.21043 PS=0.99 NRD=19.68 NRS=13.116 M=1 R=4.26667
+ SA=75001.4 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1006_d N_A_27_74#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.207307 AS=0.1036 PD=1.39957 PS=1.02 NRD=29.184 NRS=0 M=1 R=4.93333
+ SA=75001.8 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_27_74#_M1007_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 A_150_392# N_C_M1001_g N_A_27_74#_M1001_s VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1005 A_234_392# N_B_M1005_g A_150_392# VPB PSHORT L=0.15 W=1 AD=0.21 AS=0.135
+ PD=1.42 PS=1.27 NRD=30.5153 NRS=15.7403 M=1 R=6.66667 SA=75000.6 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_234_392# VPB PSHORT L=0.15 W=1 AD=0.231981
+ AS=0.21 PD=1.49057 PS=1.42 NRD=1.9503 NRS=30.5153 M=1 R=6.66667 SA=75001.2
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1002_d N_A_27_74#_M1002_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.259819 PD=1.42 PS=1.66943 NRD=1.7533 NRS=29.8849 M=1 R=7.46667
+ SA=75001.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1003 N_X_M1002_d N_A_27_74#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.1 SB=75000.3 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__or3_2.pxi.spice"
*
.ends
*
*
