* File: sky130_fd_sc_hs__sdlclkp_1.pxi.spice
* Created: Tue Sep  1 20:24:01 2020
* 
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%SCE N_SCE_c_159_n N_SCE_M1010_g N_SCE_c_164_n
+ N_SCE_M1015_g SCE N_SCE_c_161_n N_SCE_c_162_n
+ PM_SKY130_FD_SC_HS__SDLCLKP_1%SCE
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%GATE N_GATE_c_194_n N_GATE_M1005_g
+ N_GATE_M1009_g GATE N_GATE_c_196_n PM_SKY130_FD_SC_HS__SDLCLKP_1%GATE
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%A_318_74# N_A_318_74#_M1000_d
+ N_A_318_74#_M1001_d N_A_318_74#_c_241_n N_A_318_74#_M1017_g
+ N_A_318_74#_M1011_g N_A_318_74#_c_235_n N_A_318_74#_c_236_n
+ N_A_318_74#_c_237_n N_A_318_74#_c_238_n N_A_318_74#_c_239_n
+ N_A_318_74#_c_240_n PM_SKY130_FD_SC_HS__SDLCLKP_1%A_318_74#
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%A_288_48# N_A_288_48#_M1003_s
+ N_A_288_48#_M1002_s N_A_288_48#_c_311_n N_A_288_48#_M1000_g
+ N_A_288_48#_c_312_n N_A_288_48#_c_313_n N_A_288_48#_c_314_n
+ N_A_288_48#_c_331_n N_A_288_48#_c_332_n N_A_288_48#_c_333_n
+ N_A_288_48#_M1001_g N_A_288_48#_c_335_n N_A_288_48#_c_336_n
+ N_A_288_48#_c_315_n N_A_288_48#_c_316_n N_A_288_48#_c_317_n
+ N_A_288_48#_M1014_g N_A_288_48#_c_337_n N_A_288_48#_M1016_g
+ N_A_288_48#_c_338_n N_A_288_48#_c_318_n N_A_288_48#_c_319_n
+ N_A_288_48#_c_320_n N_A_288_48#_c_321_n N_A_288_48#_c_322_n
+ N_A_288_48#_c_323_n N_A_288_48#_c_379_p N_A_288_48#_c_324_n
+ N_A_288_48#_c_325_n N_A_288_48#_c_326_n N_A_288_48#_c_327_n
+ N_A_288_48#_c_328_n N_A_288_48#_c_329_n N_A_288_48#_c_340_n
+ PM_SKY130_FD_SC_HS__SDLCLKP_1%A_288_48#
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%A_709_54# N_A_709_54#_M1008_d
+ N_A_709_54#_M1012_d N_A_709_54#_M1013_g N_A_709_54#_c_493_n
+ N_A_709_54#_c_494_n N_A_709_54#_M1007_g N_A_709_54#_c_484_n
+ N_A_709_54#_M1006_g N_A_709_54#_c_485_n N_A_709_54#_c_496_n
+ N_A_709_54#_M1021_g N_A_709_54#_c_497_n N_A_709_54#_c_486_n
+ N_A_709_54#_c_487_n N_A_709_54#_c_499_n N_A_709_54#_c_500_n
+ N_A_709_54#_c_488_n N_A_709_54#_c_489_n N_A_709_54#_c_502_n
+ N_A_709_54#_c_503_n N_A_709_54#_c_490_n N_A_709_54#_c_491_n
+ N_A_709_54#_c_504_n PM_SKY130_FD_SC_HS__SDLCLKP_1%A_709_54#
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%A_566_74# N_A_566_74#_M1014_d
+ N_A_566_74#_M1017_d N_A_566_74#_c_614_n N_A_566_74#_M1008_g
+ N_A_566_74#_c_615_n N_A_566_74#_M1012_g N_A_566_74#_c_616_n
+ N_A_566_74#_c_617_n N_A_566_74#_c_618_n N_A_566_74#_c_619_n
+ N_A_566_74#_c_623_n N_A_566_74#_c_620_n
+ PM_SKY130_FD_SC_HS__SDLCLKP_1%A_566_74#
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%CLK N_CLK_M1003_g N_CLK_c_696_n N_CLK_M1002_g
+ N_CLK_M1004_g N_CLK_c_697_n N_CLK_c_694_n N_CLK_c_699_n N_CLK_M1020_g CLK
+ N_CLK_c_695_n PM_SKY130_FD_SC_HS__SDLCLKP_1%CLK
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%A_1238_94# N_A_1238_94#_M1006_d
+ N_A_1238_94#_M1020_d N_A_1238_94#_c_761_n N_A_1238_94#_M1019_g
+ N_A_1238_94#_M1018_g N_A_1238_94#_c_753_n N_A_1238_94#_c_754_n
+ N_A_1238_94#_c_755_n N_A_1238_94#_c_756_n N_A_1238_94#_c_764_n
+ N_A_1238_94#_c_757_n N_A_1238_94#_c_758_n N_A_1238_94#_c_759_n
+ N_A_1238_94#_c_760_n PM_SKY130_FD_SC_HS__SDLCLKP_1%A_1238_94#
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%VPWR N_VPWR_M1015_s N_VPWR_M1001_s
+ N_VPWR_M1007_d N_VPWR_M1002_d N_VPWR_M1021_d N_VPWR_c_819_n N_VPWR_c_820_n
+ N_VPWR_c_821_n N_VPWR_c_822_n N_VPWR_c_823_n N_VPWR_c_824_n N_VPWR_c_825_n
+ N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n VPWR N_VPWR_c_829_n
+ N_VPWR_c_830_n N_VPWR_c_831_n N_VPWR_c_818_n N_VPWR_c_833_n N_VPWR_c_834_n
+ PM_SKY130_FD_SC_HS__SDLCLKP_1%VPWR
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%A_114_112# N_A_114_112#_M1010_d
+ N_A_114_112#_M1014_s N_A_114_112#_M1005_d N_A_114_112#_M1017_s
+ N_A_114_112#_c_919_n N_A_114_112#_c_906_n N_A_114_112#_c_907_n
+ N_A_114_112#_c_908_n N_A_114_112#_c_909_n N_A_114_112#_c_910_n
+ N_A_114_112#_c_915_n N_A_114_112#_c_916_n N_A_114_112#_c_917_n
+ N_A_114_112#_c_911_n N_A_114_112#_c_918_n N_A_114_112#_c_912_n
+ N_A_114_112#_c_913_n PM_SKY130_FD_SC_HS__SDLCLKP_1%A_114_112#
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%GCLK N_GCLK_M1018_d N_GCLK_M1019_d
+ N_GCLK_c_1009_n N_GCLK_c_1010_n GCLK GCLK GCLK GCLK N_GCLK_c_1011_n
+ PM_SKY130_FD_SC_HS__SDLCLKP_1%GCLK
x_PM_SKY130_FD_SC_HS__SDLCLKP_1%VGND N_VGND_M1010_s N_VGND_M1009_d
+ N_VGND_M1013_d N_VGND_M1003_d N_VGND_M1018_s N_VGND_c_1030_n N_VGND_c_1031_n
+ N_VGND_c_1032_n N_VGND_c_1033_n N_VGND_c_1034_n N_VGND_c_1035_n
+ N_VGND_c_1036_n VGND N_VGND_c_1037_n N_VGND_c_1038_n N_VGND_c_1039_n
+ N_VGND_c_1040_n N_VGND_c_1041_n N_VGND_c_1042_n N_VGND_c_1043_n
+ N_VGND_c_1044_n PM_SKY130_FD_SC_HS__SDLCLKP_1%VGND
cc_1 VNB N_SCE_c_159_n 0.0157839f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.773
cc_2 VNB N_SCE_M1010_g 0.0259568f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_3 VNB N_SCE_c_161_n 0.0236738f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_4 VNB N_SCE_c_162_n 0.0150641f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_5 VNB N_GATE_c_194_n 0.00752289f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.477
cc_6 VNB N_GATE_M1009_g 0.0408954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_GATE_c_196_n 0.00329566f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.455
cc_8 VNB N_A_318_74#_M1011_g 0.0389156f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.455
cc_9 VNB N_A_318_74#_c_235_n 0.00339384f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.29
cc_10 VNB N_A_318_74#_c_236_n 0.00231274f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_11 VNB N_A_318_74#_c_237_n 0.00736224f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.625
cc_12 VNB N_A_318_74#_c_238_n 0.00390824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_318_74#_c_239_n 0.00408366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_318_74#_c_240_n 0.0434898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_288_48#_c_311_n 0.0220743f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_16 VNB N_A_288_48#_c_312_n 0.0226305f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_A_288_48#_c_313_n 0.00998942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_288_48#_c_314_n 0.0222673f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_19 VNB N_A_288_48#_c_315_n 0.0289975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_288_48#_c_316_n 0.0486971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_288_48#_c_317_n 0.0185017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_288_48#_c_318_n 0.00119764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_288_48#_c_319_n 0.00547716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_288_48#_c_320_n 0.00507066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_288_48#_c_321_n 3.42301e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_288_48#_c_322_n 0.00855195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_288_48#_c_323_n 0.00227124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_288_48#_c_324_n 0.0162494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_288_48#_c_325_n 0.0018167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_288_48#_c_326_n 0.00525123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_288_48#_c_327_n 0.0107853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_288_48#_c_328_n 0.0090122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_288_48#_c_329_n 0.00699471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_709_54#_M1013_g 0.0520948f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_35 VNB N_A_709_54#_c_484_n 0.0183947f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_36 VNB N_A_709_54#_c_485_n 0.00607584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_709_54#_c_486_n 0.00310352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_709_54#_c_487_n 0.00569356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_709_54#_c_488_n 0.00230943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_709_54#_c_489_n 0.00109471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_709_54#_c_490_n 0.00886798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_709_54#_c_491_n 0.0520879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_566_74#_c_614_n 0.0210688f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_44 VNB N_A_566_74#_c_615_n 0.0528587f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_45 VNB N_A_566_74#_c_616_n 0.00288593f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_46 VNB N_A_566_74#_c_617_n 0.00111963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_566_74#_c_618_n 0.0123613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_566_74#_c_619_n 0.00271082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_566_74#_c_620_n 0.00512979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_CLK_M1003_g 0.0287493f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.29
cc_51 VNB N_CLK_M1004_g 0.0225156f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_52 VNB N_CLK_c_694_n 0.0389302f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_53 VNB N_CLK_c_695_n 0.00149199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1238_94#_c_753_n 0.0203562f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_55 VNB N_A_1238_94#_c_754_n 0.0216435f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_56 VNB N_A_1238_94#_c_755_n 0.00818435f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.29
cc_57 VNB N_A_1238_94#_c_756_n 0.00126393f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_58 VNB N_A_1238_94#_c_757_n 0.00338577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1238_94#_c_758_n 0.0110227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1238_94#_c_759_n 0.0137359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1238_94#_c_760_n 0.0126688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VPWR_c_818_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_114_112#_c_906_n 0.00158689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_114_112#_c_907_n 0.00325089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_114_112#_c_908_n 0.0152342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_114_112#_c_909_n 0.00499122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_114_112#_c_910_n 0.0042758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_114_112#_c_911_n 0.00507239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_114_112#_c_912_n 0.0064939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_114_112#_c_913_n 0.00971962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_GCLK_c_1009_n 0.0264315f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_72 VNB N_GCLK_c_1010_n 0.0128764f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_73 VNB N_GCLK_c_1011_n 0.0248543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1030_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_75 VNB N_VGND_c_1031_n 0.0503666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1032_n 0.00818657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1033_n 0.0148257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1034_n 0.0138206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1035_n 0.0594191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1036_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1037_n 0.0191862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1038_n 0.0363448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1039_n 0.0336226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1040_n 0.0190343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1041_n 0.450913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1042_n 0.0174852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1043_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1044_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VPB N_SCE_c_159_n 0.0387567f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.773
cc_90 VPB N_SCE_c_164_n 0.0189667f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_91 VPB N_SCE_c_162_n 0.0123756f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_92 VPB N_GATE_c_194_n 0.0519215f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.477
cc_93 VPB N_GATE_c_196_n 0.00479274f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.455
cc_94 VPB N_A_318_74#_c_241_n 0.0177558f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_95 VPB N_A_318_74#_c_236_n 0.00391009f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.625
cc_96 VPB N_A_318_74#_c_238_n 0.0074227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_318_74#_c_239_n 0.00364869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_318_74#_c_240_n 0.0295175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_288_48#_c_314_n 9.64921e-19 $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_100 VPB N_A_288_48#_c_331_n 0.00878738f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_101 VPB N_A_288_48#_c_332_n 0.0202349f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_102 VPB N_A_288_48#_c_333_n 0.00741006f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.625
cc_103 VPB N_A_288_48#_M1001_g 0.0102552f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.625
cc_104 VPB N_A_288_48#_c_335_n 0.105598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_288_48#_c_336_n 0.0139993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_288_48#_c_337_n 0.0189875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_288_48#_c_338_n 0.0262172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_288_48#_c_327_n 0.00788597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_288_48#_c_340_n 0.00803822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_709_54#_M1013_g 0.00833695f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_111 VPB N_A_709_54#_c_493_n 0.0117917f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.455
cc_112 VPB N_A_709_54#_c_494_n 0.0211796f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_113 VPB N_A_709_54#_c_485_n 0.0111936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_709_54#_c_496_n 0.0213215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_709_54#_c_497_n 0.00621316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_709_54#_c_487_n 0.00145732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_709_54#_c_499_n 0.00422519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_709_54#_c_500_n 0.011802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_709_54#_c_488_n 0.00315495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_709_54#_c_502_n 0.00888013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_709_54#_c_503_n 0.00725981f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_709_54#_c_504_n 0.0517179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_566_74#_c_615_n 0.028466f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_124 VPB N_A_566_74#_c_617_n 0.00733186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_566_74#_c_623_n 0.00133434f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_CLK_c_696_n 0.0197057f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_127 VPB N_CLK_c_697_n 0.0216753f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.455
cc_128 VPB N_CLK_c_694_n 0.0385177f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_129 VPB N_CLK_c_699_n 0.016087f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_130 VPB N_CLK_c_695_n 0.00107524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_1238_94#_c_761_n 0.0215523f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_132 VPB N_A_1238_94#_c_755_n 0.015177f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_133 VPB N_A_1238_94#_c_756_n 0.00336531f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.625
cc_134 VPB N_A_1238_94#_c_764_n 0.00306307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_819_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.625
cc_136 VPB N_VPWR_c_820_n 0.0420655f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_821_n 0.0161505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_822_n 0.0121801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_823_n 0.0161862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_824_n 0.0105562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_825_n 0.0349499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_826_n 0.0077576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_827_n 0.0202398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_828_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_829_n 0.0312656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_830_n 0.0651369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_831_n 0.0201101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_818_n 0.105874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_833_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_834_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_114_112#_c_910_n 0.00933921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_114_112#_c_915_n 0.0134682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_114_112#_c_916_n 0.0122028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_114_112#_c_917_n 0.00644621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_114_112#_c_918_n 0.00851359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB GCLK 0.0136177f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_157 VPB GCLK 0.0416962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_GCLK_c_1011_n 0.00778299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 N_SCE_c_159_n N_GATE_c_194_n 0.0257045f $X=0.407 $Y=1.773 $X2=-0.19
+ $Y2=-0.245
cc_160 N_SCE_c_164_n N_GATE_c_194_n 0.0523559f $X=0.505 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_161 N_SCE_c_162_n N_GATE_c_194_n 0.00106303f $X=0.385 $Y=1.455 $X2=-0.19
+ $Y2=-0.245
cc_162 N_SCE_M1010_g N_GATE_M1009_g 0.0205103f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_163 N_SCE_c_161_n N_GATE_M1009_g 0.0173046f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_164 N_SCE_c_162_n N_GATE_M1009_g 0.00112397f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_165 N_SCE_c_159_n N_GATE_c_196_n 0.00179107f $X=0.407 $Y=1.773 $X2=0 $Y2=0
cc_166 N_SCE_c_164_n N_GATE_c_196_n 0.00180688f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_167 N_SCE_c_162_n N_GATE_c_196_n 0.0184673f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_168 N_SCE_c_159_n N_VPWR_c_820_n 0.00510697f $X=0.407 $Y=1.773 $X2=0 $Y2=0
cc_169 N_SCE_c_164_n N_VPWR_c_820_n 0.0214995f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_170 N_SCE_c_162_n N_VPWR_c_820_n 0.0255262f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_171 N_SCE_c_164_n N_VPWR_c_829_n 0.00413917f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_172 N_SCE_c_164_n N_VPWR_c_818_n 0.00817239f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_173 N_SCE_M1010_g N_A_114_112#_c_919_n 0.00259685f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_174 N_SCE_M1010_g N_A_114_112#_c_906_n 0.00358583f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_175 N_SCE_M1010_g N_A_114_112#_c_907_n 0.00332504f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_176 N_SCE_c_161_n N_A_114_112#_c_909_n 0.00130413f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_177 N_SCE_c_162_n N_A_114_112#_c_909_n 0.0145604f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_178 N_SCE_c_164_n N_A_114_112#_c_916_n 4.68407e-19 $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_179 N_SCE_M1010_g N_A_114_112#_c_911_n 0.00419565f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_180 N_SCE_c_161_n N_A_114_112#_c_911_n 0.00118053f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_181 N_SCE_c_164_n N_A_114_112#_c_918_n 0.00137187f $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_182 N_SCE_M1010_g N_VGND_c_1031_n 0.00819892f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_183 N_SCE_c_161_n N_VGND_c_1031_n 0.00386581f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_184 N_SCE_c_162_n N_VGND_c_1031_n 0.0216167f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_185 N_SCE_M1010_g N_VGND_c_1037_n 0.00432822f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_186 N_SCE_M1010_g N_VGND_c_1041_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_187 N_GATE_M1009_g N_A_318_74#_c_237_n 0.00108365f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_188 N_GATE_M1009_g N_A_288_48#_c_311_n 0.0251298f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_189 N_GATE_c_194_n N_VPWR_c_820_n 0.00324913f $X=0.895 $Y=2.045 $X2=0 $Y2=0
cc_190 N_GATE_c_194_n N_VPWR_c_821_n 0.00329562f $X=0.895 $Y=2.045 $X2=0 $Y2=0
cc_191 N_GATE_c_194_n N_VPWR_c_829_n 0.00445602f $X=0.895 $Y=2.045 $X2=0 $Y2=0
cc_192 N_GATE_c_194_n N_VPWR_c_818_n 0.00858051f $X=0.895 $Y=2.045 $X2=0 $Y2=0
cc_193 N_GATE_c_196_n N_A_114_112#_M1005_d 0.00267407f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_194 N_GATE_M1009_g N_A_114_112#_c_919_n 0.00510645f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_195 N_GATE_M1009_g N_A_114_112#_c_906_n 0.00455954f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_196 N_GATE_M1009_g N_A_114_112#_c_907_n 0.00216557f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_197 N_GATE_c_194_n N_A_114_112#_c_908_n 9.51679e-19 $X=0.895 $Y=2.045 $X2=0
+ $Y2=0
cc_198 N_GATE_M1009_g N_A_114_112#_c_908_n 0.009786f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_199 N_GATE_c_196_n N_A_114_112#_c_908_n 0.0314033f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_200 N_GATE_c_194_n N_A_114_112#_c_909_n 3.45023e-19 $X=0.895 $Y=2.045 $X2=0
+ $Y2=0
cc_201 N_GATE_M1009_g N_A_114_112#_c_909_n 0.00215547f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_202 N_GATE_c_196_n N_A_114_112#_c_909_n 0.00675183f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_203 N_GATE_c_194_n N_A_114_112#_c_910_n 0.00514915f $X=0.895 $Y=2.045 $X2=0
+ $Y2=0
cc_204 N_GATE_M1009_g N_A_114_112#_c_910_n 0.00428574f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_205 N_GATE_c_196_n N_A_114_112#_c_910_n 0.0424879f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_206 N_GATE_c_194_n N_A_114_112#_c_916_n 0.00361198f $X=0.895 $Y=2.045 $X2=0
+ $Y2=0
cc_207 N_GATE_c_196_n N_A_114_112#_c_916_n 0.0215997f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_208 N_GATE_M1009_g N_A_114_112#_c_911_n 0.00476476f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_209 N_GATE_c_194_n N_A_114_112#_c_918_n 0.00893078f $X=0.895 $Y=2.045 $X2=0
+ $Y2=0
cc_210 N_GATE_M1009_g N_A_114_112#_c_913_n 0.00917045f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_211 N_GATE_M1009_g N_VGND_c_1037_n 0.00340632f $X=0.925 $Y=0.835 $X2=0 $Y2=0
cc_212 N_GATE_M1009_g N_VGND_c_1041_n 0.00487769f $X=0.925 $Y=0.835 $X2=0 $Y2=0
cc_213 N_A_318_74#_c_235_n N_A_288_48#_c_311_n 0.00194041f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_214 N_A_318_74#_c_237_n N_A_288_48#_c_311_n 0.005869f $X=1.73 $Y=0.965 $X2=0
+ $Y2=0
cc_215 N_A_318_74#_c_235_n N_A_288_48#_c_312_n 0.00954194f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_216 N_A_318_74#_c_237_n N_A_288_48#_c_312_n 0.00448444f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_217 N_A_318_74#_c_238_n N_A_288_48#_c_312_n 4.8832e-19 $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_218 N_A_318_74#_c_235_n N_A_288_48#_c_314_n 0.00816401f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_219 N_A_318_74#_c_238_n N_A_288_48#_c_314_n 0.0126287f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_220 N_A_318_74#_c_239_n N_A_288_48#_c_314_n 7.2504e-19 $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_221 N_A_318_74#_c_240_n N_A_288_48#_c_314_n 0.00607965f $X=3 $Y=1.602 $X2=0
+ $Y2=0
cc_222 N_A_318_74#_c_238_n N_A_288_48#_c_333_n 0.00536326f $X=2.38 $Y=1.847
+ $X2=0 $Y2=0
cc_223 N_A_318_74#_c_238_n N_A_288_48#_M1001_g 0.0154189f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_224 N_A_318_74#_c_241_n N_A_288_48#_c_335_n 0.0103487f $X=3 $Y=1.82 $X2=0
+ $Y2=0
cc_225 N_A_318_74#_c_236_n N_A_288_48#_c_315_n 0.00115318f $X=2.625 $Y=1.63
+ $X2=0 $Y2=0
cc_226 N_A_318_74#_c_239_n N_A_288_48#_c_315_n 9.741e-19 $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_227 N_A_318_74#_c_240_n N_A_288_48#_c_315_n 0.0114346f $X=3 $Y=1.602 $X2=0
+ $Y2=0
cc_228 N_A_318_74#_c_235_n N_A_288_48#_c_316_n 0.00509279f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_229 N_A_318_74#_c_237_n N_A_288_48#_c_316_n 0.00163563f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_230 N_A_318_74#_c_238_n N_A_288_48#_c_316_n 0.0045155f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_231 N_A_318_74#_M1011_g N_A_288_48#_c_317_n 0.0224891f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_232 N_A_318_74#_c_241_n N_A_288_48#_c_337_n 0.0100718f $X=3 $Y=1.82 $X2=0
+ $Y2=0
cc_233 N_A_318_74#_M1011_g N_A_288_48#_c_318_n 0.00115934f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_234 N_A_318_74#_c_237_n N_A_288_48#_c_318_n 0.00472036f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_235 N_A_318_74#_M1011_g N_A_288_48#_c_319_n 0.0127767f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_236 N_A_318_74#_M1011_g N_A_288_48#_c_321_n 0.00543799f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_237 N_A_318_74#_M1011_g N_A_288_48#_c_323_n 0.00118267f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_238 N_A_318_74#_M1011_g N_A_288_48#_c_328_n 4.23122e-19 $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_239 N_A_318_74#_c_235_n N_A_288_48#_c_328_n 0.0176486f $X=1.88 $Y=1.545 $X2=0
+ $Y2=0
cc_240 N_A_318_74#_c_236_n N_A_288_48#_c_328_n 0.0101474f $X=2.625 $Y=1.63 $X2=0
+ $Y2=0
cc_241 N_A_318_74#_c_237_n N_A_288_48#_c_328_n 0.00760911f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_242 N_A_318_74#_c_238_n N_A_288_48#_c_328_n 0.0216474f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_243 N_A_318_74#_c_239_n N_A_288_48#_c_328_n 0.00707468f $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_244 N_A_318_74#_c_240_n N_A_288_48#_c_328_n 3.53521e-19 $X=3 $Y=1.602 $X2=0
+ $Y2=0
cc_245 N_A_318_74#_M1011_g N_A_709_54#_M1013_g 0.0878255f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_246 N_A_318_74#_c_240_n N_A_709_54#_M1013_g 0.00213846f $X=3 $Y=1.602 $X2=0
+ $Y2=0
cc_247 N_A_318_74#_c_241_n N_A_709_54#_c_504_n 0.0037268f $X=3 $Y=1.82 $X2=0
+ $Y2=0
cc_248 N_A_318_74#_M1011_g N_A_566_74#_c_616_n 0.00783189f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_249 N_A_318_74#_c_241_n N_A_566_74#_c_617_n 0.0118423f $X=3 $Y=1.82 $X2=0
+ $Y2=0
cc_250 N_A_318_74#_c_239_n N_A_566_74#_c_617_n 0.0121454f $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_251 N_A_318_74#_c_240_n N_A_566_74#_c_617_n 0.0193292f $X=3 $Y=1.602 $X2=0
+ $Y2=0
cc_252 N_A_318_74#_M1011_g N_A_566_74#_c_619_n 0.00886883f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_253 N_A_318_74#_c_239_n N_A_566_74#_c_619_n 5.28074e-19 $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_254 N_A_318_74#_c_240_n N_A_566_74#_c_619_n 0.00591219f $X=3 $Y=1.602 $X2=0
+ $Y2=0
cc_255 N_A_318_74#_c_241_n N_A_566_74#_c_623_n 0.00433065f $X=3 $Y=1.82 $X2=0
+ $Y2=0
cc_256 N_A_318_74#_M1011_g N_A_566_74#_c_620_n 0.0114381f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_257 N_A_318_74#_c_239_n N_A_566_74#_c_620_n 0.0129997f $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_258 N_A_318_74#_c_240_n N_A_566_74#_c_620_n 0.0104014f $X=3 $Y=1.602 $X2=0
+ $Y2=0
cc_259 N_A_318_74#_c_238_n N_VPWR_M1001_s 0.00401388f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_260 N_A_318_74#_c_241_n N_VPWR_c_818_n 9.39239e-19 $X=3 $Y=1.82 $X2=0 $Y2=0
cc_261 N_A_318_74#_c_235_n N_A_114_112#_c_908_n 0.0137774f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_262 N_A_318_74#_c_237_n N_A_114_112#_c_908_n 0.0048023f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_263 N_A_318_74#_c_235_n N_A_114_112#_c_910_n 0.00636232f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_264 N_A_318_74#_c_238_n N_A_114_112#_c_910_n 0.0495324f $X=2.38 $Y=1.847
+ $X2=0 $Y2=0
cc_265 N_A_318_74#_M1001_d N_A_114_112#_c_915_n 0.0056824f $X=2.065 $Y=1.84
+ $X2=0 $Y2=0
cc_266 N_A_318_74#_c_241_n N_A_114_112#_c_915_n 0.00348124f $X=3 $Y=1.82 $X2=0
+ $Y2=0
cc_267 N_A_318_74#_c_236_n N_A_114_112#_c_915_n 0.00713243f $X=2.625 $Y=1.63
+ $X2=0 $Y2=0
cc_268 N_A_318_74#_c_238_n N_A_114_112#_c_915_n 0.0370266f $X=2.38 $Y=1.847
+ $X2=0 $Y2=0
cc_269 N_A_318_74#_c_241_n N_A_114_112#_c_917_n 0.00317398f $X=3 $Y=1.82 $X2=0
+ $Y2=0
cc_270 N_A_318_74#_c_236_n N_A_114_112#_c_917_n 0.00118245f $X=2.625 $Y=1.63
+ $X2=0 $Y2=0
cc_271 N_A_318_74#_c_238_n N_A_114_112#_c_917_n 0.0182961f $X=2.38 $Y=1.847
+ $X2=0 $Y2=0
cc_272 N_A_318_74#_c_239_n N_A_114_112#_c_917_n 0.0197455f $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_273 N_A_318_74#_c_240_n N_A_114_112#_c_917_n 0.00184413f $X=3 $Y=1.602 $X2=0
+ $Y2=0
cc_274 N_A_318_74#_M1000_d N_A_114_112#_c_913_n 0.00669008f $X=1.59 $Y=0.37
+ $X2=0 $Y2=0
cc_275 N_A_318_74#_c_237_n N_A_114_112#_c_913_n 0.0255794f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_276 N_A_318_74#_M1011_g N_VGND_c_1035_n 9.29978e-19 $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_277 N_A_288_48#_c_324_n N_A_709_54#_M1008_d 0.00266942f $X=4.9 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_278 N_A_288_48#_c_319_n N_A_709_54#_M1013_g 0.00362604f $X=3.41 $Y=0.34 $X2=0
+ $Y2=0
cc_279 N_A_288_48#_c_321_n N_A_709_54#_M1013_g 0.00875253f $X=3.495 $Y=0.88
+ $X2=0 $Y2=0
cc_280 N_A_288_48#_c_322_n N_A_709_54#_M1013_g 0.0112599f $X=4.09 $Y=0.965 $X2=0
+ $Y2=0
cc_281 N_A_288_48#_c_323_n N_A_709_54#_M1013_g 0.0019606f $X=3.58 $Y=0.965 $X2=0
+ $Y2=0
cc_282 N_A_288_48#_c_379_p N_A_709_54#_M1013_g 0.00159596f $X=4.175 $Y=0.88
+ $X2=0 $Y2=0
cc_283 N_A_288_48#_c_337_n N_A_709_54#_c_494_n 0.032469f $X=3.535 $Y=2.955 $X2=0
+ $Y2=0
cc_284 N_A_288_48#_c_338_n N_A_709_54#_c_494_n 0.00318616f $X=3.535 $Y=3.15
+ $X2=0 $Y2=0
cc_285 N_A_288_48#_c_324_n N_A_709_54#_c_486_n 0.0187364f $X=4.9 $Y=0.34 $X2=0
+ $Y2=0
cc_286 N_A_288_48#_c_326_n N_A_709_54#_c_486_n 0.0181109f $X=5.065 $Y=0.515
+ $X2=0 $Y2=0
cc_287 N_A_288_48#_c_327_n N_A_709_54#_c_487_n 0.0304982f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_288 N_A_288_48#_c_340_n N_A_709_54#_c_499_n 0.0172409f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_289 N_A_288_48#_M1002_s N_A_709_54#_c_500_n 0.00789244f $X=5.07 $Y=2.015
+ $X2=0 $Y2=0
cc_290 N_A_288_48#_c_340_n N_A_709_54#_c_500_n 0.0255233f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_291 N_A_288_48#_c_327_n N_A_709_54#_c_488_n 0.00560204f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_292 N_A_288_48#_c_340_n N_A_709_54#_c_488_n 0.0115936f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_293 N_A_288_48#_c_329_n N_A_709_54#_c_489_n 0.0181109f $X=5.065 $Y=1.13 $X2=0
+ $Y2=0
cc_294 N_A_288_48#_c_327_n N_A_709_54#_c_502_n 0.0215371f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_295 N_A_288_48#_c_340_n N_A_709_54#_c_502_n 0.0111525f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_296 N_A_288_48#_c_327_n N_A_709_54#_c_490_n 0.00357445f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_297 N_A_288_48#_c_337_n N_A_709_54#_c_504_n 0.00535945f $X=3.535 $Y=2.955
+ $X2=0 $Y2=0
cc_298 N_A_288_48#_c_319_n N_A_566_74#_M1014_d 0.00256812f $X=3.41 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_299 N_A_288_48#_c_322_n N_A_566_74#_c_614_n 0.00554178f $X=4.09 $Y=0.965
+ $X2=0 $Y2=0
cc_300 N_A_288_48#_c_379_p N_A_566_74#_c_614_n 0.0123114f $X=4.175 $Y=0.88 $X2=0
+ $Y2=0
cc_301 N_A_288_48#_c_324_n N_A_566_74#_c_614_n 0.0114613f $X=4.9 $Y=0.34 $X2=0
+ $Y2=0
cc_302 N_A_288_48#_c_325_n N_A_566_74#_c_614_n 0.00278978f $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_303 N_A_288_48#_c_326_n N_A_566_74#_c_614_n 0.00362229f $X=5.065 $Y=0.515
+ $X2=0 $Y2=0
cc_304 N_A_288_48#_c_322_n N_A_566_74#_c_615_n 0.00521109f $X=4.09 $Y=0.965
+ $X2=0 $Y2=0
cc_305 N_A_288_48#_c_327_n N_A_566_74#_c_615_n 0.00200979f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_306 N_A_288_48#_c_340_n N_A_566_74#_c_615_n 5.53173e-19 $X=5.215 $Y=2.16
+ $X2=0 $Y2=0
cc_307 N_A_288_48#_c_316_n N_A_566_74#_c_616_n 2.9126e-19 $X=2.415 $Y=1.07 $X2=0
+ $Y2=0
cc_308 N_A_288_48#_c_317_n N_A_566_74#_c_616_n 0.00183864f $X=2.755 $Y=0.995
+ $X2=0 $Y2=0
cc_309 N_A_288_48#_c_318_n N_A_566_74#_c_616_n 0.00430473f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_310 N_A_288_48#_c_323_n N_A_566_74#_c_616_n 0.0100841f $X=3.58 $Y=0.965 $X2=0
+ $Y2=0
cc_311 N_A_288_48#_c_328_n N_A_566_74#_c_616_n 0.00848118f $X=2.25 $Y=1.195
+ $X2=0 $Y2=0
cc_312 N_A_288_48#_c_337_n N_A_566_74#_c_617_n 0.00760144f $X=3.535 $Y=2.955
+ $X2=0 $Y2=0
cc_313 N_A_288_48#_c_322_n N_A_566_74#_c_618_n 0.0502793f $X=4.09 $Y=0.965 $X2=0
+ $Y2=0
cc_314 N_A_288_48#_c_323_n N_A_566_74#_c_618_n 0.0147362f $X=3.58 $Y=0.965 $X2=0
+ $Y2=0
cc_315 N_A_288_48#_c_318_n N_A_566_74#_c_619_n 0.0112956f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_316 N_A_288_48#_c_319_n N_A_566_74#_c_619_n 0.0209617f $X=3.41 $Y=0.34 $X2=0
+ $Y2=0
cc_317 N_A_288_48#_c_321_n N_A_566_74#_c_619_n 0.021236f $X=3.495 $Y=0.88 $X2=0
+ $Y2=0
cc_318 N_A_288_48#_c_323_n N_A_566_74#_c_619_n 0.00374694f $X=3.58 $Y=0.965
+ $X2=0 $Y2=0
cc_319 N_A_288_48#_c_335_n N_A_566_74#_c_623_n 0.0064175f $X=3.445 $Y=3.15 $X2=0
+ $Y2=0
cc_320 N_A_288_48#_c_316_n N_A_566_74#_c_620_n 8.48984e-19 $X=2.415 $Y=1.07
+ $X2=0 $Y2=0
cc_321 N_A_288_48#_c_328_n N_A_566_74#_c_620_n 0.00421113f $X=2.25 $Y=1.195
+ $X2=0 $Y2=0
cc_322 N_A_288_48#_c_324_n N_CLK_M1003_g 0.0047004f $X=4.9 $Y=0.34 $X2=0 $Y2=0
cc_323 N_A_288_48#_c_326_n N_CLK_M1003_g 0.00681907f $X=5.065 $Y=0.515 $X2=0
+ $Y2=0
cc_324 N_A_288_48#_c_327_n N_CLK_M1003_g 0.0109213f $X=5.075 $Y=1.995 $X2=0
+ $Y2=0
cc_325 N_A_288_48#_c_329_n N_CLK_M1003_g 0.00328501f $X=5.065 $Y=1.13 $X2=0
+ $Y2=0
cc_326 N_A_288_48#_c_327_n N_CLK_c_696_n 0.00124615f $X=5.075 $Y=1.995 $X2=0
+ $Y2=0
cc_327 N_A_288_48#_c_340_n N_CLK_c_696_n 0.00616665f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_328 N_A_288_48#_c_327_n N_CLK_c_694_n 0.00549078f $X=5.075 $Y=1.995 $X2=0
+ $Y2=0
cc_329 N_A_288_48#_c_340_n N_CLK_c_694_n 0.00539247f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_330 N_A_288_48#_c_327_n N_CLK_c_695_n 0.0323289f $X=5.075 $Y=1.995 $X2=0
+ $Y2=0
cc_331 N_A_288_48#_c_340_n N_CLK_c_695_n 0.00334638f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_332 N_A_288_48#_c_331_n N_VPWR_c_821_n 0.0195176f $X=1.99 $Y=2.845 $X2=0
+ $Y2=0
cc_333 N_A_288_48#_M1001_g N_VPWR_c_821_n 0.00391084f $X=1.99 $Y=2.26 $X2=0
+ $Y2=0
cc_334 N_A_288_48#_c_337_n N_VPWR_c_822_n 0.00188736f $X=3.535 $Y=2.955 $X2=0
+ $Y2=0
cc_335 N_A_288_48#_c_338_n N_VPWR_c_822_n 0.00576281f $X=3.535 $Y=3.15 $X2=0
+ $Y2=0
cc_336 N_A_288_48#_c_336_n N_VPWR_c_830_n 0.0555583f $X=2.08 $Y=3.15 $X2=0 $Y2=0
cc_337 N_A_288_48#_c_335_n N_VPWR_c_818_n 0.0415959f $X=3.445 $Y=3.15 $X2=0
+ $Y2=0
cc_338 N_A_288_48#_c_336_n N_VPWR_c_818_n 0.00793983f $X=2.08 $Y=3.15 $X2=0
+ $Y2=0
cc_339 N_A_288_48#_c_338_n N_VPWR_c_818_n 0.0132593f $X=3.535 $Y=3.15 $X2=0
+ $Y2=0
cc_340 N_A_288_48#_c_318_n N_A_114_112#_M1014_s 0.0084363f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_341 N_A_288_48#_c_320_n N_A_114_112#_M1014_s 6.08643e-19 $X=2.715 $Y=0.34
+ $X2=0 $Y2=0
cc_342 N_A_288_48#_c_311_n N_A_114_112#_c_919_n 0.00137149f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_343 N_A_288_48#_c_312_n N_A_114_112#_c_908_n 0.00258488f $X=1.9 $Y=1.285
+ $X2=0 $Y2=0
cc_344 N_A_288_48#_c_313_n N_A_114_112#_c_908_n 0.00935869f $X=1.59 $Y=1.285
+ $X2=0 $Y2=0
cc_345 N_A_288_48#_c_314_n N_A_114_112#_c_908_n 6.11401e-19 $X=1.99 $Y=1.675
+ $X2=0 $Y2=0
cc_346 N_A_288_48#_c_314_n N_A_114_112#_c_910_n 0.00164805f $X=1.99 $Y=1.675
+ $X2=0 $Y2=0
cc_347 N_A_288_48#_M1001_g N_A_114_112#_c_910_n 0.00717054f $X=1.99 $Y=2.26
+ $X2=0 $Y2=0
cc_348 N_A_288_48#_M1001_g N_A_114_112#_c_915_n 0.0225531f $X=1.99 $Y=2.26 $X2=0
+ $Y2=0
cc_349 N_A_288_48#_c_335_n N_A_114_112#_c_915_n 0.0163697f $X=3.445 $Y=3.15
+ $X2=0 $Y2=0
cc_350 N_A_288_48#_M1001_g N_A_114_112#_c_917_n 0.00377738f $X=1.99 $Y=2.26
+ $X2=0 $Y2=0
cc_351 N_A_288_48#_c_313_n N_A_114_112#_c_911_n 0.00137149f $X=1.59 $Y=1.285
+ $X2=0 $Y2=0
cc_352 N_A_288_48#_M1001_g N_A_114_112#_c_918_n 0.00405881f $X=1.99 $Y=2.26
+ $X2=0 $Y2=0
cc_353 N_A_288_48#_c_311_n N_A_114_112#_c_912_n 0.00622457f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_354 N_A_288_48#_c_316_n N_A_114_112#_c_912_n 0.00597962f $X=2.415 $Y=1.07
+ $X2=0 $Y2=0
cc_355 N_A_288_48#_c_317_n N_A_114_112#_c_912_n 0.00235306f $X=2.755 $Y=0.995
+ $X2=0 $Y2=0
cc_356 N_A_288_48#_c_318_n N_A_114_112#_c_912_n 0.0276253f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_357 N_A_288_48#_c_320_n N_A_114_112#_c_912_n 0.00627272f $X=2.715 $Y=0.34
+ $X2=0 $Y2=0
cc_358 N_A_288_48#_c_328_n N_A_114_112#_c_912_n 0.0142183f $X=2.25 $Y=1.195
+ $X2=0 $Y2=0
cc_359 N_A_288_48#_c_311_n N_A_114_112#_c_913_n 0.0154871f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_360 N_A_288_48#_c_312_n N_A_114_112#_c_913_n 7.62669e-19 $X=1.9 $Y=1.285
+ $X2=0 $Y2=0
cc_361 N_A_288_48#_c_316_n N_A_114_112#_c_913_n 0.00222971f $X=2.415 $Y=1.07
+ $X2=0 $Y2=0
cc_362 N_A_288_48#_c_322_n N_VGND_M1013_d 0.00663756f $X=4.09 $Y=0.965 $X2=0
+ $Y2=0
cc_363 N_A_288_48#_c_379_p N_VGND_M1013_d 0.00488787f $X=4.175 $Y=0.88 $X2=0
+ $Y2=0
cc_364 N_A_288_48#_c_325_n N_VGND_M1013_d 5.22721e-19 $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_365 N_A_288_48#_c_319_n N_VGND_c_1032_n 0.01267f $X=3.41 $Y=0.34 $X2=0 $Y2=0
cc_366 N_A_288_48#_c_322_n N_VGND_c_1032_n 0.013847f $X=4.09 $Y=0.965 $X2=0
+ $Y2=0
cc_367 N_A_288_48#_c_379_p N_VGND_c_1032_n 0.020664f $X=4.175 $Y=0.88 $X2=0
+ $Y2=0
cc_368 N_A_288_48#_c_325_n N_VGND_c_1032_n 0.0142265f $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_369 N_A_288_48#_c_324_n N_VGND_c_1033_n 0.0112234f $X=4.9 $Y=0.34 $X2=0 $Y2=0
cc_370 N_A_288_48#_c_326_n N_VGND_c_1033_n 0.0259244f $X=5.065 $Y=0.515 $X2=0
+ $Y2=0
cc_371 N_A_288_48#_c_311_n N_VGND_c_1035_n 0.00315544f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_372 N_A_288_48#_c_317_n N_VGND_c_1035_n 0.00278237f $X=2.755 $Y=0.995 $X2=0
+ $Y2=0
cc_373 N_A_288_48#_c_319_n N_VGND_c_1035_n 0.0565673f $X=3.41 $Y=0.34 $X2=0
+ $Y2=0
cc_374 N_A_288_48#_c_320_n N_VGND_c_1035_n 0.0120637f $X=2.715 $Y=0.34 $X2=0
+ $Y2=0
cc_375 N_A_288_48#_c_324_n N_VGND_c_1038_n 0.0644063f $X=4.9 $Y=0.34 $X2=0 $Y2=0
cc_376 N_A_288_48#_c_325_n N_VGND_c_1038_n 0.0120637f $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_377 N_A_288_48#_c_311_n N_VGND_c_1041_n 0.00400711f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_378 N_A_288_48#_c_317_n N_VGND_c_1041_n 0.00363424f $X=2.755 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_288_48#_c_319_n N_VGND_c_1041_n 0.0322089f $X=3.41 $Y=0.34 $X2=0
+ $Y2=0
cc_380 N_A_288_48#_c_320_n N_VGND_c_1041_n 0.00644906f $X=2.715 $Y=0.34 $X2=0
+ $Y2=0
cc_381 N_A_288_48#_c_324_n N_VGND_c_1041_n 0.036247f $X=4.9 $Y=0.34 $X2=0 $Y2=0
cc_382 N_A_288_48#_c_325_n N_VGND_c_1041_n 0.00644906f $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_383 N_A_288_48#_c_311_n N_VGND_c_1042_n 0.00542971f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_384 N_A_288_48#_c_319_n A_667_80# 6.48644e-19 $X=3.41 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_385 N_A_288_48#_c_321_n A_667_80# 0.00370274f $X=3.495 $Y=0.88 $X2=-0.19
+ $Y2=-0.245
cc_386 N_A_709_54#_M1013_g N_A_566_74#_c_614_n 0.0149957f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_387 N_A_709_54#_c_487_n N_A_566_74#_c_614_n 0.00622278f $X=4.585 $Y=1.74
+ $X2=0 $Y2=0
cc_388 N_A_709_54#_M1013_g N_A_566_74#_c_615_n 0.0190415f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_389 N_A_709_54#_c_494_n N_A_566_74#_c_615_n 0.0119201f $X=3.925 $Y=2.385
+ $X2=0 $Y2=0
cc_390 N_A_709_54#_c_497_n N_A_566_74#_c_615_n 0.0320047f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_391 N_A_709_54#_c_487_n N_A_566_74#_c_615_n 0.0216923f $X=4.585 $Y=1.74 $X2=0
+ $Y2=0
cc_392 N_A_709_54#_c_499_n N_A_566_74#_c_615_n 0.006408f $X=4.655 $Y=2.495 $X2=0
+ $Y2=0
cc_393 N_A_709_54#_c_489_n N_A_566_74#_c_615_n 0.00269107f $X=4.555 $Y=1.05
+ $X2=0 $Y2=0
cc_394 N_A_709_54#_c_502_n N_A_566_74#_c_615_n 0.00129855f $X=4.655 $Y=1.905
+ $X2=0 $Y2=0
cc_395 N_A_709_54#_c_503_n N_A_566_74#_c_615_n 0.00497499f $X=4.655 $Y=2.58
+ $X2=0 $Y2=0
cc_396 N_A_709_54#_c_504_n N_A_566_74#_c_615_n 0.0229405f $X=3.925 $Y=1.955
+ $X2=0 $Y2=0
cc_397 N_A_709_54#_M1013_g N_A_566_74#_c_616_n 0.00101991f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_398 N_A_709_54#_M1013_g N_A_566_74#_c_617_n 0.00820694f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_399 N_A_709_54#_c_493_n N_A_566_74#_c_617_n 0.00598811f $X=3.925 $Y=2.295
+ $X2=0 $Y2=0
cc_400 N_A_709_54#_c_497_n N_A_566_74#_c_617_n 0.0269421f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_401 N_A_709_54#_M1013_g N_A_566_74#_c_618_n 0.0175999f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_402 N_A_709_54#_c_497_n N_A_566_74#_c_618_n 0.0538499f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_403 N_A_709_54#_c_487_n N_A_566_74#_c_618_n 0.0251783f $X=4.585 $Y=1.74 $X2=0
+ $Y2=0
cc_404 N_A_709_54#_c_504_n N_A_566_74#_c_618_n 0.00190817f $X=3.925 $Y=1.955
+ $X2=0 $Y2=0
cc_405 N_A_709_54#_M1013_g N_A_566_74#_c_619_n 2.77632e-19 $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_406 N_A_709_54#_c_486_n N_CLK_M1003_g 0.00101752f $X=4.515 $Y=0.82 $X2=0
+ $Y2=0
cc_407 N_A_709_54#_c_490_n N_CLK_M1003_g 3.97134e-19 $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_408 N_A_709_54#_c_499_n N_CLK_c_696_n 0.00394589f $X=4.655 $Y=2.495 $X2=0
+ $Y2=0
cc_409 N_A_709_54#_c_500_n N_CLK_c_696_n 0.0185052f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_410 N_A_709_54#_c_488_n N_CLK_c_696_n 0.00665398f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_411 N_A_709_54#_c_502_n N_CLK_c_696_n 3.42277e-19 $X=4.655 $Y=1.905 $X2=0
+ $Y2=0
cc_412 N_A_709_54#_c_503_n N_CLK_c_696_n 0.00628162f $X=4.655 $Y=2.58 $X2=0
+ $Y2=0
cc_413 N_A_709_54#_c_484_n N_CLK_M1004_g 0.0365055f $X=6.115 $Y=1.22 $X2=0 $Y2=0
cc_414 N_A_709_54#_c_490_n N_CLK_M1004_g 0.00389357f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_415 N_A_709_54#_c_485_n N_CLK_c_697_n 0.00711822f $X=6.585 $Y=1.85 $X2=0
+ $Y2=0
cc_416 N_A_709_54#_c_488_n N_CLK_c_697_n 0.0148834f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_417 N_A_709_54#_c_490_n N_CLK_c_697_n 0.00356342f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_418 N_A_709_54#_c_491_n N_CLK_c_697_n 0.0117835f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_419 N_A_709_54#_c_485_n N_CLK_c_694_n 0.0025851f $X=6.585 $Y=1.85 $X2=0 $Y2=0
cc_420 N_A_709_54#_c_500_n N_CLK_c_694_n 0.00623917f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_421 N_A_709_54#_c_488_n N_CLK_c_694_n 0.00388892f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_422 N_A_709_54#_c_491_n N_CLK_c_694_n 0.0365055f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_423 N_A_709_54#_c_496_n N_CLK_c_699_n 0.0147207f $X=6.585 $Y=1.94 $X2=0 $Y2=0
cc_424 N_A_709_54#_c_500_n N_CLK_c_699_n 0.00197375f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_425 N_A_709_54#_c_488_n N_CLK_c_699_n 0.00575084f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_426 N_A_709_54#_c_488_n N_CLK_c_695_n 0.0172833f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_427 N_A_709_54#_c_490_n N_CLK_c_695_n 0.0150518f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_428 N_A_709_54#_c_485_n N_A_1238_94#_c_761_n 0.00596996f $X=6.585 $Y=1.85
+ $X2=0 $Y2=0
cc_429 N_A_709_54#_c_496_n N_A_1238_94#_c_761_n 0.0175258f $X=6.585 $Y=1.94
+ $X2=0 $Y2=0
cc_430 N_A_709_54#_c_491_n N_A_1238_94#_c_753_n 0.00914688f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_431 N_A_709_54#_c_485_n N_A_1238_94#_c_755_n 0.0105675f $X=6.585 $Y=1.85
+ $X2=0 $Y2=0
cc_432 N_A_709_54#_c_485_n N_A_1238_94#_c_756_n 0.0108131f $X=6.585 $Y=1.85
+ $X2=0 $Y2=0
cc_433 N_A_709_54#_c_496_n N_A_1238_94#_c_756_n 0.00780012f $X=6.585 $Y=1.94
+ $X2=0 $Y2=0
cc_434 N_A_709_54#_c_488_n N_A_1238_94#_c_756_n 0.0184253f $X=5.915 $Y=2.495
+ $X2=0 $Y2=0
cc_435 N_A_709_54#_c_490_n N_A_1238_94#_c_756_n 0.0297948f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_436 N_A_709_54#_c_491_n N_A_1238_94#_c_756_n 0.0163379f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_437 N_A_709_54#_c_496_n N_A_1238_94#_c_764_n 0.0152265f $X=6.585 $Y=1.94
+ $X2=0 $Y2=0
cc_438 N_A_709_54#_c_500_n N_A_1238_94#_c_764_n 0.0126254f $X=5.83 $Y=2.58 $X2=0
+ $Y2=0
cc_439 N_A_709_54#_c_488_n N_A_1238_94#_c_764_n 0.0400627f $X=5.915 $Y=2.495
+ $X2=0 $Y2=0
cc_440 N_A_709_54#_c_484_n N_A_1238_94#_c_757_n 0.00421972f $X=6.115 $Y=1.22
+ $X2=0 $Y2=0
cc_441 N_A_709_54#_c_490_n N_A_1238_94#_c_757_n 0.00580698f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_442 N_A_709_54#_c_491_n N_A_1238_94#_c_757_n 0.00749726f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_443 N_A_709_54#_c_485_n N_A_1238_94#_c_758_n 0.0023274f $X=6.585 $Y=1.85
+ $X2=0 $Y2=0
cc_444 N_A_709_54#_c_491_n N_A_1238_94#_c_758_n 0.00244172f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_445 N_A_709_54#_c_491_n N_A_1238_94#_c_759_n 0.00899294f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_446 N_A_709_54#_c_484_n N_A_1238_94#_c_760_n 0.0110552f $X=6.115 $Y=1.22
+ $X2=0 $Y2=0
cc_447 N_A_709_54#_c_490_n N_A_1238_94#_c_760_n 0.00874612f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_448 N_A_709_54#_c_491_n N_A_1238_94#_c_760_n 0.0075575f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_449 N_A_709_54#_c_497_n N_VPWR_M1007_d 0.00304656f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_450 N_A_709_54#_c_500_n N_VPWR_M1002_d 0.0138319f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_451 N_A_709_54#_c_488_n N_VPWR_M1002_d 0.0139379f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_452 N_A_709_54#_c_494_n N_VPWR_c_822_n 0.0131507f $X=3.925 $Y=2.385 $X2=0
+ $Y2=0
cc_453 N_A_709_54#_c_497_n N_VPWR_c_822_n 0.0170087f $X=4.49 $Y=1.93 $X2=0 $Y2=0
cc_454 N_A_709_54#_c_499_n N_VPWR_c_822_n 0.0176013f $X=4.655 $Y=2.495 $X2=0
+ $Y2=0
cc_455 N_A_709_54#_c_500_n N_VPWR_c_823_n 0.0322115f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_456 N_A_709_54#_c_496_n N_VPWR_c_824_n 0.00762087f $X=6.585 $Y=1.94 $X2=0
+ $Y2=0
cc_457 N_A_709_54#_c_500_n N_VPWR_c_825_n 0.0116981f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_458 N_A_709_54#_c_503_n N_VPWR_c_825_n 0.0110196f $X=4.655 $Y=2.58 $X2=0
+ $Y2=0
cc_459 N_A_709_54#_c_496_n N_VPWR_c_827_n 0.00491343f $X=6.585 $Y=1.94 $X2=0
+ $Y2=0
cc_460 N_A_709_54#_c_494_n N_VPWR_c_830_n 0.00467292f $X=3.925 $Y=2.385 $X2=0
+ $Y2=0
cc_461 N_A_709_54#_c_494_n N_VPWR_c_818_n 0.00471987f $X=3.925 $Y=2.385 $X2=0
+ $Y2=0
cc_462 N_A_709_54#_c_496_n N_VPWR_c_818_n 0.00512916f $X=6.585 $Y=1.94 $X2=0
+ $Y2=0
cc_463 N_A_709_54#_c_500_n N_VPWR_c_818_n 0.0233651f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_464 N_A_709_54#_c_503_n N_VPWR_c_818_n 0.0114996f $X=4.655 $Y=2.58 $X2=0
+ $Y2=0
cc_465 N_A_709_54#_M1013_g N_VGND_c_1032_n 0.0012897f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_466 N_A_709_54#_c_484_n N_VGND_c_1034_n 0.00313422f $X=6.115 $Y=1.22 $X2=0
+ $Y2=0
cc_467 N_A_709_54#_M1013_g N_VGND_c_1035_n 0.00447942f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_468 N_A_709_54#_c_484_n N_VGND_c_1039_n 0.00485498f $X=6.115 $Y=1.22 $X2=0
+ $Y2=0
cc_469 N_A_709_54#_M1013_g N_VGND_c_1041_n 0.0041113f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_470 N_A_709_54#_c_484_n N_VGND_c_1041_n 0.00514438f $X=6.115 $Y=1.22 $X2=0
+ $Y2=0
cc_471 N_A_566_74#_c_615_n N_CLK_M1003_g 0.00465657f $X=4.43 $Y=1.685 $X2=0
+ $Y2=0
cc_472 N_A_566_74#_c_615_n N_VPWR_c_822_n 0.0056644f $X=4.43 $Y=1.685 $X2=0
+ $Y2=0
cc_473 N_A_566_74#_c_623_n N_VPWR_c_822_n 0.00913742f $X=3.225 $Y=2.59 $X2=0
+ $Y2=0
cc_474 N_A_566_74#_c_615_n N_VPWR_c_825_n 0.00507376f $X=4.43 $Y=1.685 $X2=0
+ $Y2=0
cc_475 N_A_566_74#_c_623_n N_VPWR_c_830_n 0.00731246f $X=3.225 $Y=2.59 $X2=0
+ $Y2=0
cc_476 N_A_566_74#_c_615_n N_VPWR_c_818_n 0.00520574f $X=4.43 $Y=1.685 $X2=0
+ $Y2=0
cc_477 N_A_566_74#_c_623_n N_VPWR_c_818_n 0.00906972f $X=3.225 $Y=2.59 $X2=0
+ $Y2=0
cc_478 N_A_566_74#_c_617_n N_A_114_112#_c_915_n 0.00731865f $X=3.225 $Y=2.05
+ $X2=0 $Y2=0
cc_479 N_A_566_74#_c_623_n N_A_114_112#_c_915_n 0.0226116f $X=3.225 $Y=2.59
+ $X2=0 $Y2=0
cc_480 N_A_566_74#_c_617_n N_A_114_112#_c_917_n 0.0280129f $X=3.225 $Y=2.05
+ $X2=0 $Y2=0
cc_481 N_A_566_74#_c_614_n N_VGND_c_1032_n 0.00168945f $X=4.3 $Y=1.22 $X2=0
+ $Y2=0
cc_482 N_A_566_74#_c_614_n N_VGND_c_1038_n 0.00278237f $X=4.3 $Y=1.22 $X2=0
+ $Y2=0
cc_483 N_A_566_74#_c_614_n N_VGND_c_1041_n 0.00363424f $X=4.3 $Y=1.22 $X2=0
+ $Y2=0
cc_484 N_CLK_c_697_n N_A_1238_94#_c_756_n 0.00309887f $X=6.06 $Y=1.865 $X2=0
+ $Y2=0
cc_485 N_CLK_c_696_n N_A_1238_94#_c_764_n 9.17516e-19 $X=5.44 $Y=1.94 $X2=0
+ $Y2=0
cc_486 N_CLK_c_697_n N_A_1238_94#_c_764_n 0.00180466f $X=6.06 $Y=1.865 $X2=0
+ $Y2=0
cc_487 N_CLK_c_699_n N_A_1238_94#_c_764_n 0.0148784f $X=6.135 $Y=1.94 $X2=0
+ $Y2=0
cc_488 N_CLK_M1004_g N_A_1238_94#_c_760_n 0.00166928f $X=5.755 $Y=0.79 $X2=0
+ $Y2=0
cc_489 N_CLK_c_696_n N_VPWR_c_823_n 0.00460974f $X=5.44 $Y=1.94 $X2=0 $Y2=0
cc_490 N_CLK_c_699_n N_VPWR_c_823_n 0.00382137f $X=6.135 $Y=1.94 $X2=0 $Y2=0
cc_491 N_CLK_c_696_n N_VPWR_c_825_n 0.00389135f $X=5.44 $Y=1.94 $X2=0 $Y2=0
cc_492 N_CLK_c_699_n N_VPWR_c_827_n 0.00491343f $X=6.135 $Y=1.94 $X2=0 $Y2=0
cc_493 N_CLK_c_696_n N_VPWR_c_818_n 0.00512916f $X=5.44 $Y=1.94 $X2=0 $Y2=0
cc_494 N_CLK_c_699_n N_VPWR_c_818_n 0.00512916f $X=6.135 $Y=1.94 $X2=0 $Y2=0
cc_495 N_CLK_M1003_g N_VGND_c_1033_n 0.00310756f $X=5.28 $Y=0.74 $X2=0 $Y2=0
cc_496 N_CLK_M1004_g N_VGND_c_1033_n 0.00381172f $X=5.755 $Y=0.79 $X2=0 $Y2=0
cc_497 N_CLK_c_694_n N_VGND_c_1033_n 0.00109716f $X=5.83 $Y=1.865 $X2=0 $Y2=0
cc_498 N_CLK_c_695_n N_VGND_c_1033_n 0.0173191f $X=5.495 $Y=1.52 $X2=0 $Y2=0
cc_499 N_CLK_M1003_g N_VGND_c_1038_n 0.00430908f $X=5.28 $Y=0.74 $X2=0 $Y2=0
cc_500 N_CLK_M1004_g N_VGND_c_1039_n 0.00507111f $X=5.755 $Y=0.79 $X2=0 $Y2=0
cc_501 N_CLK_M1003_g N_VGND_c_1041_n 0.0082568f $X=5.28 $Y=0.74 $X2=0 $Y2=0
cc_502 N_CLK_M1004_g N_VGND_c_1041_n 0.00514438f $X=5.755 $Y=0.79 $X2=0 $Y2=0
cc_503 N_A_1238_94#_c_764_n N_VPWR_c_823_n 0.00276433f $X=6.36 $Y=2.16 $X2=0
+ $Y2=0
cc_504 N_A_1238_94#_c_761_n N_VPWR_c_824_n 0.0190358f $X=7.09 $Y=1.765 $X2=0
+ $Y2=0
cc_505 N_A_1238_94#_c_755_n N_VPWR_c_824_n 0.00183643f $X=7.09 $Y=1.55 $X2=0
+ $Y2=0
cc_506 N_A_1238_94#_c_764_n N_VPWR_c_824_n 0.0313712f $X=6.36 $Y=2.16 $X2=0
+ $Y2=0
cc_507 N_A_1238_94#_c_758_n N_VPWR_c_824_n 0.0123479f $X=7.08 $Y=1.465 $X2=0
+ $Y2=0
cc_508 N_A_1238_94#_c_764_n N_VPWR_c_827_n 0.0101887f $X=6.36 $Y=2.16 $X2=0
+ $Y2=0
cc_509 N_A_1238_94#_c_761_n N_VPWR_c_831_n 0.00429299f $X=7.09 $Y=1.765 $X2=0
+ $Y2=0
cc_510 N_A_1238_94#_c_761_n N_VPWR_c_818_n 0.00851465f $X=7.09 $Y=1.765 $X2=0
+ $Y2=0
cc_511 N_A_1238_94#_c_764_n N_VPWR_c_818_n 0.0112927f $X=6.36 $Y=2.16 $X2=0
+ $Y2=0
cc_512 N_A_1238_94#_c_754_n N_GCLK_c_1009_n 0.00840121f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_513 N_A_1238_94#_c_754_n N_GCLK_c_1010_n 0.00343235f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_514 N_A_1238_94#_c_761_n GCLK 0.0299017f $X=7.09 $Y=1.765 $X2=0 $Y2=0
cc_515 N_A_1238_94#_c_755_n GCLK 0.00132156f $X=7.09 $Y=1.55 $X2=0 $Y2=0
cc_516 N_A_1238_94#_c_756_n GCLK 0.00211506f $X=6.36 $Y=1.89 $X2=0 $Y2=0
cc_517 N_A_1238_94#_c_758_n GCLK 6.98006e-19 $X=7.08 $Y=1.465 $X2=0 $Y2=0
cc_518 N_A_1238_94#_c_754_n N_GCLK_c_1011_n 0.0159294f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_519 N_A_1238_94#_c_755_n N_GCLK_c_1011_n 0.00130385f $X=7.09 $Y=1.55 $X2=0
+ $Y2=0
cc_520 N_A_1238_94#_c_758_n N_GCLK_c_1011_n 0.0261275f $X=7.08 $Y=1.465 $X2=0
+ $Y2=0
cc_521 N_A_1238_94#_c_760_n N_VGND_c_1033_n 0.0101545f $X=6.33 $Y=0.615 $X2=0
+ $Y2=0
cc_522 N_A_1238_94#_c_753_n N_VGND_c_1034_n 0.00449375f $X=7.09 $Y=1.36 $X2=0
+ $Y2=0
cc_523 N_A_1238_94#_c_754_n N_VGND_c_1034_n 0.0196053f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_524 N_A_1238_94#_c_758_n N_VGND_c_1034_n 0.0213215f $X=7.08 $Y=1.465 $X2=0
+ $Y2=0
cc_525 N_A_1238_94#_c_760_n N_VGND_c_1034_n 0.0556027f $X=6.33 $Y=0.615 $X2=0
+ $Y2=0
cc_526 N_A_1238_94#_c_760_n N_VGND_c_1039_n 0.0150236f $X=6.33 $Y=0.615 $X2=0
+ $Y2=0
cc_527 N_A_1238_94#_c_754_n N_VGND_c_1040_n 0.00434272f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_528 N_A_1238_94#_c_754_n N_VGND_c_1041_n 0.00828811f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_529 N_A_1238_94#_c_760_n N_VGND_c_1041_n 0.0164774f $X=6.33 $Y=0.615 $X2=0
+ $Y2=0
cc_530 N_VPWR_M1001_s N_A_114_112#_c_910_n 0.00750857f $X=1.535 $Y=1.84 $X2=0
+ $Y2=0
cc_531 N_VPWR_M1001_s N_A_114_112#_c_915_n 0.0107006f $X=1.535 $Y=1.84 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_830_n N_A_114_112#_c_915_n 0.00575553f $X=3.985 $Y=3.33 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_818_n N_A_114_112#_c_915_n 0.0301793f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_534 N_VPWR_M1001_s N_A_114_112#_c_916_n 0.00203332f $X=1.535 $Y=1.84 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_820_n N_A_114_112#_c_916_n 0.0054501f $X=0.28 $Y=2.295 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_821_n N_A_114_112#_c_916_n 0.0260892f $X=1.68 $Y=2.825 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_818_n N_A_114_112#_c_916_n 0.00909594f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_820_n N_A_114_112#_c_918_n 0.0149893f $X=0.28 $Y=2.295 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_821_n N_A_114_112#_c_918_n 0.0215742f $X=1.68 $Y=2.825 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_829_n N_A_114_112#_c_918_n 0.0142535f $X=1.515 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_818_n N_A_114_112#_c_918_n 0.0119151f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_824_n GCLK 0.0610124f $X=6.86 $Y=2.225 $X2=0 $Y2=0
cc_543 N_VPWR_c_831_n GCLK 0.0155281f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_544 N_VPWR_c_818_n GCLK 0.0128528f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_545 N_A_114_112#_c_913_n N_VGND_M1009_d 0.00979382f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_546 N_A_114_112#_c_919_n N_VGND_c_1031_n 0.0150351f $X=0.71 $Y=0.83 $X2=0
+ $Y2=0
cc_547 N_A_114_112#_c_907_n N_VGND_c_1031_n 0.00756924f $X=0.885 $Y=0.625 $X2=0
+ $Y2=0
cc_548 N_A_114_112#_c_912_n N_VGND_c_1035_n 0.0107474f $X=2.29 $Y=0.565 $X2=0
+ $Y2=0
cc_549 N_A_114_112#_c_913_n N_VGND_c_1035_n 0.0151341f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_550 N_A_114_112#_c_907_n N_VGND_c_1037_n 0.0083132f $X=0.885 $Y=0.625 $X2=0
+ $Y2=0
cc_551 N_A_114_112#_c_913_n N_VGND_c_1037_n 0.00360867f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_552 N_A_114_112#_c_907_n N_VGND_c_1041_n 0.0109521f $X=0.885 $Y=0.625 $X2=0
+ $Y2=0
cc_553 N_A_114_112#_c_912_n N_VGND_c_1041_n 0.00908767f $X=2.29 $Y=0.565 $X2=0
+ $Y2=0
cc_554 N_A_114_112#_c_913_n N_VGND_c_1041_n 0.0289707f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_555 N_A_114_112#_c_913_n N_VGND_c_1042_n 0.0242087f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_556 N_GCLK_c_1009_n N_VGND_c_1034_n 0.0302381f $X=7.405 $Y=0.515 $X2=0 $Y2=0
cc_557 N_GCLK_c_1009_n N_VGND_c_1040_n 0.0152332f $X=7.405 $Y=0.515 $X2=0 $Y2=0
cc_558 N_GCLK_c_1009_n N_VGND_c_1041_n 0.0125524f $X=7.405 $Y=0.515 $X2=0 $Y2=0
