* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nor2b_1 A B_N VGND VNB VPB VPWR Y
M1000 VPWR B_N a_27_112# VPB pshort w=840000u l=150000u
+  ad=4.69e+11p pd=3.16e+06u as=2.478e+11p ps=2.27e+06u
M1001 a_278_368# A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1002 VGND a_27_112# Y VNB nlowvt w=740000u l=150000u
+  ad=5.6985e+11p pd=4.59e+06u as=2.627e+11p ps=2.19e+06u
M1003 VGND B_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.805e+11p ps=2.12e+06u
M1004 Y a_27_112# a_278_368# VPB pshort w=1.12e+06u l=150000u
+  ad=4.2e+11p pd=2.99e+06u as=0p ps=0u
M1005 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
