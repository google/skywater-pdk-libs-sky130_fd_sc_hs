* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__and3b_4 A_N B C VGND VNB VPB VPWR X
X0 a_298_368# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_239_98# B a_498_98# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 X a_298_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 X a_298_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 a_298_368# a_27_74# a_239_98# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 VPWR B a_298_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 a_298_368# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 VGND C a_498_98# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VPWR C a_298_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X9 VPWR a_298_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X10 VPWR a_298_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X11 a_498_98# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 VGND a_298_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_298_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X14 VPWR a_27_74# a_298_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X15 VGND a_298_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_498_98# B a_239_98# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X18 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_239_98# a_27_74# a_298_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 X a_298_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 X a_298_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
