* File: sky130_fd_sc_hs__dlxbn_1.pex.spice
* Created: Tue Sep  1 20:02:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DLXBN_1%D 3 5 6 8 9 12 14
c37 6 0 2.98693e-19 $X=0.675 $Y=2.045
r38 12 14 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.592 $Y=1.425
+ $X2=0.592 $Y2=1.26
r39 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6
+ $Y=1.425 $X2=0.6 $Y2=1.425
r40 9 13 2.14223 $w=6.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.595 $X2=0.6
+ $Y2=1.595
r41 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.675 $Y=2.045
+ $X2=0.675 $Y2=2.54
r42 5 6 49.7604 $w=2.78e-07 $l=3.25868e-07 $layer=POLY_cond $X=0.592 $Y=1.758
+ $X2=0.675 $Y2=2.045
r43 4 12 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=0.592 $Y=1.432
+ $X2=0.592 $Y2=1.425
r44 4 5 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=0.592 $Y=1.432
+ $X2=0.592 $Y2=1.758
r45 3 14 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.495 $Y=0.875
+ $X2=0.495 $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%GATE_N 3 5 7 8 12
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.795 $X2=1.17 $Y2=1.795
r37 8 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.17 $Y=2.035 $X2=1.17
+ $Y2=1.795
r38 5 11 52.2586 $w=2.99e-07 $l=2.52488e-07 $layer=POLY_cond $X=1.175 $Y=2.045
+ $X2=1.17 $Y2=1.795
r39 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.175 $Y=2.045
+ $X2=1.175 $Y2=2.54
r40 1 11 38.5562 $w=2.99e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.085 $Y=1.63
+ $X2=1.17 $Y2=1.795
r41 1 3 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.085 $Y=1.63
+ $X2=1.085 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%A_232_82# 1 2 7 9 11 13 14 16 17 19 20 21 23
+ 24 26 27 30 36 39 44 48 49 50 56 58
c131 48 0 1.69272e-19 $X=1.4 $Y=2.405
c132 17 0 1.82525e-19 $X=3.19 $Y=1.11
c133 7 0 1.72289e-19 $X=2.145 $Y=1.325
r134 53 56 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.94 $Y=1.635
+ $X2=4.06 $Y2=1.635
r135 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.635 $X2=3.94 $Y2=1.635
r136 48 50 1.83343 $w=4.38e-07 $l=7e-08 $layer=LI1_cond $X=1.455 $Y=2.405
+ $X2=1.455 $Y2=2.475
r137 48 49 6.73996 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=2.405
+ $X2=1.455 $Y2=2.32
r138 45 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.74 $Y=1.415
+ $X2=1.74 $Y2=1.325
r139 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.415 $X2=1.74 $Y2=1.415
r140 42 44 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.59 $Y=1.39
+ $X2=1.74 $Y2=1.39
r141 38 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=1.8
+ $X2=4.06 $Y2=1.635
r142 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.06 $Y=1.8 $X2=4.06
+ $Y2=2.39
r143 37 50 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.675 $Y=2.475
+ $X2=1.455 $Y2=2.475
r144 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.975 $Y=2.475
+ $X2=4.06 $Y2=2.39
r145 36 37 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.975 $Y=2.475
+ $X2=1.675 $Y2=2.475
r146 34 42 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.59 $Y=1.52
+ $X2=1.59 $Y2=1.39
r147 34 49 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.59 $Y=1.52 $X2=1.59
+ $Y2=2.32
r148 28 42 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.3 $Y=1.39
+ $X2=1.59 $Y2=1.39
r149 28 30 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.3 $Y=1.26
+ $X2=1.3 $Y2=1.005
r150 24 54 50.653 $w=3.43e-07 $l=2.68328e-07 $layer=POLY_cond $X=3.95 $Y=1.885
+ $X2=3.912 $Y2=1.635
r151 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.95 $Y=1.885
+ $X2=3.95 $Y2=2.17
r152 23 54 38.7084 $w=3.43e-07 $l=2.15708e-07 $layer=POLY_cond $X=3.795 $Y=1.47
+ $X2=3.912 $Y2=1.635
r153 22 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.795 $Y=1.26
+ $X2=3.795 $Y2=1.47
r154 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.72 $Y=1.185
+ $X2=3.795 $Y2=1.26
r155 20 21 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.72 $Y=1.185
+ $X2=3.265 $Y2=1.185
r156 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.19 $Y=1.11
+ $X2=3.265 $Y2=1.185
r157 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.19 $Y=1.11
+ $X2=3.19 $Y2=0.715
r158 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.235 $Y=1.885
+ $X2=2.235 $Y2=2.38
r159 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.235 $Y=1.795
+ $X2=2.235 $Y2=1.885
r160 12 27 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.235 $Y=1.4
+ $X2=2.235 $Y2=1.325
r161 12 13 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.235 $Y=1.4
+ $X2=2.235 $Y2=1.795
r162 9 27 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.22 $Y=1.25
+ $X2=2.235 $Y2=1.325
r163 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.22 $Y=1.25 $X2=2.22
+ $Y2=0.77
r164 8 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.325
+ $X2=1.74 $Y2=1.325
r165 7 27 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.145 $Y=1.325
+ $X2=2.235 $Y2=1.325
r166 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.145 $Y=1.325
+ $X2=1.905 $Y2=1.325
r167 2 48 300 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=2 $X=1.25
+ $Y=2.12 $X2=1.4 $Y2=2.405
r168 1 30 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.41 $X2=1.3 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%A_27_120# 1 2 8 9 11 14 20 24 25 27 33 34
c78 34 0 1.29422e-19 $X=0.32 $Y=2.1
c79 24 0 4.43268e-20 $X=2.7 $Y=1.415
c80 20 0 3.54814e-19 $X=2.535 $Y=0.665
c81 14 0 3.06626e-19 $X=2.8 $Y=0.715
c82 9 0 1.66542e-19 $X=2.78 $Y=1.885
r83 33 34 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=2.265
+ $X2=0.32 $Y2=2.1
r84 31 34 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.18 $Y=1.09
+ $X2=0.18 $Y2=2.1
r85 30 31 11.4519 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.27 $Y=0.835
+ $X2=0.27 $Y2=1.09
r86 27 30 5.59758 $w=3.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.27 $Y=0.665
+ $X2=0.27 $Y2=0.835
r87 25 37 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.415
+ $X2=2.705 $Y2=1.58
r88 25 36 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.415
+ $X2=2.705 $Y2=1.25
r89 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.415 $X2=2.7 $Y2=1.415
r90 22 24 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=2.7 $Y=0.75 $X2=2.7
+ $Y2=1.415
r91 21 27 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=0.665
+ $X2=0.27 $Y2=0.665
r92 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.535 $Y=0.665
+ $X2=2.7 $Y2=0.75
r93 20 21 136.353 $w=1.68e-07 $l=2.09e-06 $layer=LI1_cond $X=2.535 $Y=0.665
+ $X2=0.445 $Y2=0.665
r94 14 36 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.8 $Y=0.715 $X2=2.8
+ $Y2=1.25
r95 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.78 $Y=1.885
+ $X2=2.78 $Y2=2.46
r96 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.78 $Y=1.795 $X2=2.78
+ $Y2=1.885
r97 8 37 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=2.78 $Y=1.795
+ $X2=2.78 $Y2=1.58
r98 2 33 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=0.25
+ $Y=2.12 $X2=0.38 $Y2=2.265
r99 1 30 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.6 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%A_343_80# 1 2 7 9 12 13 18 19 20 22 23 25 26
+ 31 38
c98 25 0 6.89381e-20 $X=4.095 $Y=0.34
c99 18 0 1.48832e-19 $X=2.16 $Y=1.71
c100 13 0 1.57795e-19 $X=2.075 $Y=1.005
c101 7 0 4.43268e-20 $X=3.2 $Y=1.885
r102 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.635 $X2=3.25 $Y2=1.635
r103 31 33 3.93548 $w=4.03e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.845
+ $X2=3.25 $Y2=1.845
r104 29 30 4.44175 $w=4.12e-07 $l=1.5e-07 $layer=LI1_cond $X=2.01 $Y=1.965
+ $X2=2.16 $Y2=1.965
r105 26 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=0.34
+ $X2=4.095 $Y2=0.505
r106 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.095
+ $Y=0.34 $X2=4.095 $Y2=0.34
r107 23 25 41.027 $w=2.48e-07 $l=8.9e-07 $layer=LI1_cond $X=3.205 $Y=0.38
+ $X2=4.095 $Y2=0.38
r108 22 31 5.82385 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=3.12 $Y=1.47
+ $X2=3.12 $Y2=1.845
r109 21 23 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.12 $Y=0.505
+ $X2=3.205 $Y2=0.38
r110 21 22 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=3.12 $Y=0.505
+ $X2=3.12 $Y2=1.47
r111 20 30 2.51946 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=1.965
+ $X2=2.16 $Y2=1.965
r112 19 31 11.6947 $w=5.1e-07 $l=5.2156e-07 $layer=LI1_cond $X=2.655 $Y=1.965
+ $X2=3.12 $Y2=1.845
r113 19 20 9.61553 $w=5.08e-07 $l=4.1e-07 $layer=LI1_cond $X=2.655 $Y=1.965
+ $X2=2.245 $Y2=1.965
r114 18 30 5.95845 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.16 $Y=1.71
+ $X2=2.16 $Y2=1.965
r115 17 18 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.16 $Y=1.09
+ $X2=2.16 $Y2=1.71
r116 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.075 $Y=1.005
+ $X2=2.16 $Y2=1.09
r117 13 15 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.075 $Y=1.005
+ $X2=1.93 $Y2=1.005
r118 12 38 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.185 $Y=0.825
+ $X2=4.185 $Y2=0.505
r119 7 34 52.2586 $w=2.99e-07 $l=2.73861e-07 $layer=POLY_cond $X=3.2 $Y=1.885
+ $X2=3.25 $Y2=1.635
r120 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.2 $Y=1.885 $X2=3.2
+ $Y2=2.46
r121 2 29 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.96 $X2=2.01 $Y2=2.12
r122 1 15 182 $w=1.7e-07 $l=7.04344e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.4 $X2=1.93 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%A_863_294# 1 2 7 9 12 14 16 17 19 20 21 22
+ 24 25 27 28 33 37 39 41 46 48 53
c116 48 0 5.45732e-20 $X=4.48 $Y=1.635
c117 12 0 6.89381e-20 $X=4.575 $Y=0.825
r118 55 57 13.3156 $w=3.39e-07 $l=3.7e-07 $layer=LI1_cond $X=5.505 $Y=1.435
+ $X2=5.505 $Y2=1.805
r119 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.625
+ $Y=1.435 $X2=5.625 $Y2=1.435
r120 48 51 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.48 $Y=1.635
+ $X2=4.48 $Y2=1.805
r121 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.48
+ $Y=1.635 $X2=4.48 $Y2=1.635
r122 46 55 8.96717 $w=3.39e-07 $l=1.79374e-07 $layer=LI1_cond $X=5.475 $Y=1.27
+ $X2=5.505 $Y2=1.435
r123 46 53 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.475 $Y=1.27
+ $X2=5.475 $Y2=0.96
r124 41 43 28.1332 $w=3.38e-07 $l=8.3e-07 $layer=LI1_cond $X=5.39 $Y=1.905
+ $X2=5.39 $Y2=2.735
r125 39 57 3.05 $w=3.4e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.39 $Y=1.89
+ $X2=5.505 $Y2=1.805
r126 39 41 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=5.39 $Y=1.89
+ $X2=5.39 $Y2=1.905
r127 35 53 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=5.382 $Y=0.783
+ $X2=5.382 $Y2=0.96
r128 35 37 8.05087 $w=3.53e-07 $l=2.48e-07 $layer=LI1_cond $X=5.382 $Y=0.783
+ $X2=5.382 $Y2=0.535
r129 34 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=1.805
+ $X2=4.48 $Y2=1.805
r130 33 57 4.78362 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=5.22 $Y=1.805
+ $X2=5.505 $Y2=1.805
r131 33 34 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.22 $Y=1.805
+ $X2=4.645 $Y2=1.805
r132 29 30 1.59956 $w=4.52e-07 $l=1.5e-08 $layer=POLY_cond $X=6.155 $Y=1.475
+ $X2=6.17 $Y2=1.475
r133 28 56 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=6.065 $Y=1.435
+ $X2=5.625 $Y2=1.435
r134 28 29 13.1977 $w=4.52e-07 $l=1.08167e-07 $layer=POLY_cond $X=6.065 $Y=1.435
+ $X2=6.155 $Y2=1.475
r135 25 32 28.877 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.68 $Y=1.185
+ $X2=6.68 $Y2=1.475
r136 25 27 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.68 $Y=1.185
+ $X2=6.68 $Y2=0.835
r137 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.66 $Y=2.045
+ $X2=6.66 $Y2=2.54
r138 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.66 $Y=1.955
+ $X2=6.66 $Y2=2.045
r139 20 32 2.13274 $w=4.52e-07 $l=2e-08 $layer=POLY_cond $X=6.66 $Y=1.475
+ $X2=6.68 $Y2=1.475
r140 20 30 52.2522 $w=4.52e-07 $l=4.9e-07 $layer=POLY_cond $X=6.66 $Y=1.475
+ $X2=6.17 $Y2=1.475
r141 20 21 137.992 $w=1.8e-07 $l=3.55e-07 $layer=POLY_cond $X=6.66 $Y=1.6
+ $X2=6.66 $Y2=1.955
r142 17 30 28.877 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.17 $Y=1.185
+ $X2=6.17 $Y2=1.475
r143 17 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.17 $Y=1.185
+ $X2=6.17 $Y2=0.74
r144 14 29 28.877 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.155 $Y=1.765
+ $X2=6.155 $Y2=1.475
r145 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.155 $Y=1.765
+ $X2=6.155 $Y2=2.4
r146 10 49 38.5416 $w=3.03e-07 $l=2.06325e-07 $layer=POLY_cond $X=4.575 $Y=1.47
+ $X2=4.482 $Y2=1.635
r147 10 12 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.575 $Y=1.47
+ $X2=4.575 $Y2=0.825
r148 7 49 52.063 $w=3.03e-07 $l=2.72489e-07 $layer=POLY_cond $X=4.435 $Y=1.885
+ $X2=4.482 $Y2=1.635
r149 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.435 $Y=1.885
+ $X2=4.435 $Y2=2.17
r150 2 43 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.76 $X2=5.385 $Y2=2.735
r151 2 41 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.76 $X2=5.385 $Y2=1.905
r152 1 37 91 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.37 $X2=5.37 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%A_653_79# 1 2 7 9 10 12 14 15 16 18 22
c70 18 0 1.66542e-19 $X=3.53 $Y=2.135
c71 14 0 5.45732e-20 $X=3.595 $Y=2.05
r72 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.055
+ $Y=1.385 $X2=5.055 $Y2=1.385
r73 22 25 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.055 $Y=1.215
+ $X2=5.055 $Y2=1.385
r74 19 21 8.61582 $w=5.31e-07 $l=3.75e-07 $layer=LI1_cond $X=3.595 $Y=1.012
+ $X2=3.97 $Y2=1.012
r75 16 21 9.90492 $w=5.31e-07 $l=2.7332e-07 $layer=LI1_cond $X=4.135 $Y=1.215
+ $X2=3.97 $Y2=1.012
r76 15 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.89 $Y=1.215
+ $X2=5.055 $Y2=1.215
r77 15 16 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.89 $Y=1.215
+ $X2=4.135 $Y2=1.215
r78 14 18 0.716491 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.595 $Y=2.05
+ $X2=3.53 $Y2=2.135
r79 13 19 7.53601 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=3.595 $Y=1.3
+ $X2=3.595 $Y2=1.012
r80 13 14 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.595 $Y=1.3
+ $X2=3.595 $Y2=2.05
r81 10 26 59.7291 $w=3.07e-07 $l=3.42053e-07 $layer=POLY_cond $X=5.16 $Y=1.685
+ $X2=5.07 $Y2=1.385
r82 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.16 $Y=1.685
+ $X2=5.16 $Y2=2.32
r83 7 26 38.5336 $w=3.07e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.145 $Y=1.22
+ $X2=5.07 $Y2=1.385
r84 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.145 $Y=1.22 $X2=5.145
+ $Y2=0.74
r85 2 18 600 $w=1.7e-07 $l=3.31134e-07 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=1.96 $X2=3.53 $Y2=2.135
r86 1 21 91 $w=1.7e-07 $l=9.19783e-07 $layer=licon1_NDIFF $count=2 $X=3.265
+ $Y=0.395 $X2=3.97 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%A_1347_424# 1 2 7 9 12 15 19 23 27 30
r46 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.335
+ $Y=1.465 $X2=7.335 $Y2=1.465
r47 25 30 1.47678 $w=3.3e-07 $l=1.73e-07 $layer=LI1_cond $X=7.065 $Y=1.465
+ $X2=6.892 $Y2=1.465
r48 25 27 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.065 $Y=1.465
+ $X2=7.335 $Y2=1.465
r49 21 30 5.00808 $w=3.42e-07 $l=1.65e-07 $layer=LI1_cond $X=6.892 $Y=1.63
+ $X2=6.892 $Y2=1.465
r50 21 23 21.2116 $w=3.43e-07 $l=6.35e-07 $layer=LI1_cond $X=6.892 $Y=1.63
+ $X2=6.892 $Y2=2.265
r51 17 30 5.00808 $w=3.42e-07 $l=1.65997e-07 $layer=LI1_cond $X=6.89 $Y=1.3
+ $X2=6.892 $Y2=1.465
r52 17 19 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=6.89 $Y=1.3
+ $X2=6.89 $Y2=0.835
r53 15 28 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=7.565 $Y=1.465
+ $X2=7.335 $Y2=1.465
r54 15 16 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.465
+ $X2=7.655 $Y2=1.3
r55 12 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.67 $Y=0.74
+ $X2=7.67 $Y2=1.3
r56 7 15 118.763 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=7.655 $Y=1.765
+ $X2=7.655 $Y2=1.465
r57 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.655 $Y=1.765
+ $X2=7.655 $Y2=2.4
r58 2 23 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=6.735
+ $Y=2.12 $X2=6.89 $Y2=2.265
r59 1 19 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=6.755
+ $Y=0.56 $X2=6.895 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%VPWR 1 2 3 4 5 18 22 24 28 34 38 43 44 46 47
+ 49 50 51 57 75 76 79 82
r85 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r88 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r89 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r90 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r91 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r92 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r93 67 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r95 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r96 64 82 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=5.02 $Y=3.33 $X2=4.75
+ $Y2=3.33
r97 64 66 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=5.02 $Y=3.33 $X2=5.04
+ $Y2=3.33
r98 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r100 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r102 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 57 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.545 $Y2=3.33
r104 57 62 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 55 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r106 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 51 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r108 51 80 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 49 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=6.96 $Y2=3.33
r110 49 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.39 $Y2=3.33
r111 48 75 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.92 $Y2=3.33
r112 48 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.39 $Y2=3.33
r113 46 69 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.3 $Y=3.33 $X2=6
+ $Y2=3.33
r114 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.3 $Y=3.33
+ $X2=6.425 $Y2=3.33
r115 45 72 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.55 $Y=3.33
+ $X2=6.96 $Y2=3.33
r116 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.55 $Y=3.33
+ $X2=6.425 $Y2=3.33
r117 43 54 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.9 $Y2=3.33
r119 42 59 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.9 $Y2=3.33
r121 38 41 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.39 $Y=1.985
+ $X2=7.39 $Y2=2.815
r122 36 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.39 $Y=3.245
+ $X2=7.39 $Y2=3.33
r123 36 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.39 $Y=3.245
+ $X2=7.39 $Y2=2.815
r124 32 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=3.245
+ $X2=6.425 $Y2=3.33
r125 32 34 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=6.425 $Y=3.245
+ $X2=6.425 $Y2=2.265
r126 28 31 12.4038 $w=5.38e-07 $l=5.6e-07 $layer=LI1_cond $X=4.75 $Y=2.175
+ $X2=4.75 $Y2=2.735
r127 26 82 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=3.245
+ $X2=4.75 $Y2=3.33
r128 26 31 11.2963 $w=5.38e-07 $l=5.1e-07 $layer=LI1_cond $X=4.75 $Y=3.245
+ $X2=4.75 $Y2=2.735
r129 25 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.545 $Y2=3.33
r130 24 82 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=4.48 $Y=3.33
+ $X2=4.75 $Y2=3.33
r131 24 25 115.476 $w=1.68e-07 $l=1.77e-06 $layer=LI1_cond $X=4.48 $Y=3.33
+ $X2=2.71 $Y2=3.33
r132 20 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.33
r133 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=2.815
r134 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=3.245 $X2=0.9
+ $Y2=3.33
r135 16 18 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=0.9 $Y=3.245
+ $X2=0.9 $Y2=2.405
r136 5 41 400 $w=1.7e-07 $l=1.03797e-06 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.84 $X2=7.43 $Y2=2.815
r137 5 38 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.84 $X2=7.43 $Y2=1.985
r138 4 34 300 $w=1.7e-07 $l=4.96488e-07 $layer=licon1_PDIFF $count=2 $X=6.23
+ $Y=1.84 $X2=6.385 $Y2=2.265
r139 3 31 600 $w=1.7e-07 $l=9.64365e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.96 $X2=4.935 $Y2=2.735
r140 3 28 600 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.96 $X2=4.75 $Y2=2.175
r141 2 22 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=1.96 $X2=2.545 $Y2=2.815
r142 1 18 300 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=2 $X=0.75
+ $Y=2.12 $X2=0.9 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%Q 1 2 9 14 15 16 17 28
r38 21 28 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=5.96 $Y=0.93 $X2=5.96
+ $Y2=0.925
r39 17 30 7.28558 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=5.96 $Y=0.97
+ $X2=5.96 $Y2=1.1
r40 17 21 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=5.96 $Y=0.97 $X2=5.96
+ $Y2=0.93
r41 17 28 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=5.96 $Y=0.885 $X2=5.96
+ $Y2=0.925
r42 16 17 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=5.96 $Y=0.515
+ $X2=5.96 $Y2=0.885
r43 15 30 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.045 $Y=1.82
+ $X2=6.045 $Y2=1.1
r44 14 15 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.947 $Y=1.985
+ $X2=5.947 $Y2=1.82
r45 7 14 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=5.947 $Y=2.002
+ $X2=5.947 $Y2=1.985
r46 7 9 25.6695 $w=3.63e-07 $l=8.13e-07 $layer=LI1_cond $X=5.947 $Y=2.002
+ $X2=5.947 $Y2=2.815
r47 2 14 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.84 $X2=5.93 $Y2=1.985
r48 2 9 400 $w=1.7e-07 $l=1.03797e-06 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.84 $X2=5.93 $Y2=2.815
r49 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.81
+ $Y=0.37 $X2=5.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%Q_N 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=2.405
+ $X2=7.882 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.882 $Y=1.985
+ $X2=7.882 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=7.882 $Y=1.665
+ $X2=7.882 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=1.295
+ $X2=7.882 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=0.925
+ $X2=7.882 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=7.882 $Y=0.515
+ $X2=7.882 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.84 $X2=7.88 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.84 $X2=7.88 $Y2=1.985
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.745
+ $Y=0.37 $X2=7.885 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLXBN_1%VGND 1 2 3 4 5 18 22 26 29 30 32 33 34 36 41
+ 59 65 66 70 83
r79 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r80 70 73 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.79
+ $Y2=0.325
r81 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r82 66 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r83 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r84 63 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.54 $Y=0 $X2=7.415
+ $Y2=0
r85 63 65 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.54 $Y=0 $X2=7.92
+ $Y2=0
r86 62 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r87 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 59 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=7.415
+ $Y2=0
r89 59 61 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=6.96
+ $Y2=0
r90 58 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r91 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r92 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r93 54 57 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6 $Y2=0
r94 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r95 52 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r96 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r97 49 51 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=2.675 $Y=0
+ $X2=4.56 $Y2=0
r98 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r99 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r100 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r101 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r102 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r103 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r104 42 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r105 42 44 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r106 41 80 11.1804 $w=3.33e-07 $l=3.25e-07 $layer=LI1_cond $X=2.507 $Y=0
+ $X2=2.507 $Y2=0.325
r107 41 49 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.507 $Y=0
+ $X2=2.675 $Y2=0
r108 41 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r109 41 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.16
+ $Y2=0
r110 39 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r111 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r112 36 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r113 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r114 34 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r115 34 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r116 32 57 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.3 $Y=0 $X2=6 $Y2=0
r117 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.3 $Y=0 $X2=6.425
+ $Y2=0
r118 31 61 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.55 $Y=0 $X2=6.96
+ $Y2=0
r119 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.55 $Y=0 $X2=6.425
+ $Y2=0
r120 29 51 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=0
+ $X2=4.56 $Y2=0
r121 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.87
+ $Y2=0
r122 28 54 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.04
+ $Y2=0
r123 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=4.87
+ $Y2=0
r124 24 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=0.085
+ $X2=7.415 $Y2=0
r125 24 26 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.415 $Y=0.085
+ $X2=7.415 $Y2=0.515
r126 20 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=0.085
+ $X2=6.425 $Y2=0
r127 20 22 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=6.425 $Y=0.085
+ $X2=6.425 $Y2=0.89
r128 16 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0
r129 16 18 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0.535
r130 5 26 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.31
+ $Y=0.37 $X2=7.455 $Y2=0.515
r131 4 22 182 $w=1.7e-07 $l=6.05475e-07 $layer=licon1_NDIFF $count=1 $X=6.245
+ $Y=0.37 $X2=6.43 $Y2=0.89
r132 3 18 91 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=2 $X=4.65
+ $Y=0.615 $X2=4.87 $Y2=0.535
r133 2 80 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.4 $X2=2.505 $Y2=0.325
r134 1 73 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.6 $X2=0.79 $Y2=0.325
.ends

