* File: sky130_fd_sc_hs__sdfxbp_2.pex.spice
* Created: Tue Sep  1 20:23:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_36_74# 1 2 9 11 13 14 16 19 22 23 24 28
+ 36 39
c84 39 0 9.34686e-20 $X=2.03 $Y=1.89
c85 36 0 3.1124e-19 $X=0.83 $Y=1.635
c86 14 0 1.92539e-19 $X=0.965 $Y=1.635
r87 39 42 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=1.89
+ $X2=2.03 $Y2=2.055
r88 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.89 $X2=2.03 $Y2=1.89
r89 34 36 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.75 $Y=1.635 $X2=0.83
+ $Y2=1.635
r90 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.635 $X2=0.75 $Y2=1.635
r91 25 28 4.70075 $w=3.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.17 $Y=0.54
+ $X2=0.325 $Y2=0.54
r92 23 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=2.055
+ $X2=2.03 $Y2=2.055
r93 23 24 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=1.865 $Y=2.055
+ $X2=0.915 $Y2=2.055
r94 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.83 $Y=1.97
+ $X2=0.915 $Y2=2.055
r95 21 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.83 $Y=1.8 $X2=0.83
+ $Y2=1.635
r96 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.83 $Y=1.8 $X2=0.83
+ $Y2=1.97
r97 17 34 15.6453 $w=3.28e-07 $l=4.48e-07 $layer=LI1_cond $X=0.302 $Y=1.635
+ $X2=0.75 $Y2=1.635
r98 17 30 4.60977 $w=3.28e-07 $l=1.32e-07 $layer=LI1_cond $X=0.302 $Y=1.635
+ $X2=0.17 $Y2=1.635
r99 17 19 16.1607 $w=4.33e-07 $l=6.1e-07 $layer=LI1_cond $X=0.302 $Y=1.8
+ $X2=0.302 $Y2=2.41
r100 16 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=1.47
+ $X2=0.17 $Y2=1.635
r101 15 25 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.17 $Y=0.73
+ $X2=0.17 $Y2=0.54
r102 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.17 $Y=0.73
+ $X2=0.17 $Y2=1.47
r103 14 35 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.635
+ $X2=0.75 $Y2=1.635
r104 11 40 61.4066 $w=2.86e-07 $l=3.04959e-07 $layer=POLY_cond $X=2.04 $Y=2.19
+ $X2=2.03 $Y2=1.89
r105 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.04 $Y=2.19
+ $X2=2.04 $Y2=2.585
r106 7 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.04 $Y=1.47
+ $X2=0.965 $Y2=1.635
r107 7 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.04 $Y=1.47 $X2=1.04
+ $Y2=0.58
r108 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.21
+ $Y=2.265 $X2=0.355 $Y2=2.41
r109 1 28 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.37 $X2=0.325 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%SCE 2 3 4 5 7 8 10 11 13 15 16 18 19 20 24
+ 26 30 38
c75 11 0 1.11484e-19 $X=1.04 $Y=2.115
r76 32 34 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.27 $Y=1.065
+ $X2=0.54 $Y2=1.065
r77 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.065 $X2=1.91 $Y2=1.065
r78 26 30 6.311 $w=4.18e-07 $l=2.3e-07 $layer=LI1_cond $X=1.68 $Y=1.02 $X2=1.91
+ $Y2=1.02
r79 26 38 3.71646 $w=4.18e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.02
+ $X2=1.565 $Y2=1.02
r80 24 34 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.59 $Y=1.065 $X2=0.54
+ $Y2=1.065
r81 23 38 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=0.59 $Y=1.065
+ $X2=1.565 $Y2=1.065
r82 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.065 $X2=0.59 $Y2=1.065
r83 20 29 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.1 $Y=1.065
+ $X2=1.91 $Y2=1.065
r84 16 20 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.175 $Y=0.9
+ $X2=2.1 $Y2=1.065
r85 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.175 $Y=0.9
+ $X2=2.175 $Y2=0.58
r86 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.115 $Y=2.19
+ $X2=1.115 $Y2=2.585
r87 12 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.74 $Y=2.115
+ $X2=0.665 $Y2=2.115
r88 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.04 $Y=2.115
+ $X2=1.115 $Y2=2.19
r89 11 12 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.04 $Y=2.115 $X2=0.74
+ $Y2=2.115
r90 8 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.665 $Y=2.19
+ $X2=0.665 $Y2=2.115
r91 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.665 $Y=2.19
+ $X2=0.665 $Y2=2.585
r92 5 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=0.9 $X2=0.54
+ $Y2=1.065
r93 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.9 $X2=0.54
+ $Y2=0.58
r94 3 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.59 $Y=2.115
+ $X2=0.665 $Y2=2.115
r95 3 4 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.59 $Y=2.115
+ $X2=0.345 $Y2=2.115
r96 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.27 $Y=2.04
+ $X2=0.345 $Y2=2.115
r97 1 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.23
+ $X2=0.27 $Y2=1.065
r98 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.27 $Y=1.23 $X2=0.27
+ $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%D 3 6 7 9 10 13 14
c41 13 0 2.93225e-19 $X=1.49 $Y=1.635
r42 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.635
+ $X2=1.49 $Y2=1.8
r43 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.635
+ $X2=1.49 $Y2=1.47
r44 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.635 $X2=1.49 $Y2=1.635
r45 10 14 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.635
+ $X2=1.49 $Y2=1.635
r46 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.535 $Y=2.19
+ $X2=1.535 $Y2=2.585
r47 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.535 $Y=2.1 $X2=1.535
+ $Y2=2.19
r48 6 16 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=1.535 $Y=2.1 $X2=1.535
+ $Y2=1.8
r49 3 15 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.43 $Y=0.58 $X2=1.43
+ $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%SCD 1 3 6 8 12
c33 6 0 2.59705e-19 $X=2.565 $Y=0.58
c34 1 0 6.78066e-20 $X=2.525 $Y=2.19
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.94 $X2=2.57 $Y2=1.94
r36 8 12 3.12806 $w=3.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=2.035
+ $X2=2.58 $Y2=1.94
r37 4 11 38.5562 $w=2.99e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.565 $Y=1.775
+ $X2=2.57 $Y2=1.94
r38 4 6 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=2.565 $Y=1.775
+ $X2=2.565 $Y2=0.58
r39 1 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.525 $Y=2.19
+ $X2=2.57 $Y2=1.94
r40 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.525 $Y=2.19
+ $X2=2.525 $Y2=2.585
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%CLK 3 5 7 8 11
c37 11 0 6.34765e-20 $X=3.235 $Y=1.557
c38 8 0 1.30658e-19 $X=3.6 $Y=1.665
c39 5 0 1.29047e-19 $X=3.235 $Y=1.765
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.515 $X2=3.43 $Y2=1.515
r41 11 13 30.2219 $w=3.11e-07 $l=1.95e-07 $layer=POLY_cond $X=3.235 $Y=1.557
+ $X2=3.43 $Y2=1.557
r42 8 14 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.43
+ $Y2=1.565
r43 5 11 19.8172 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.235 $Y=1.765
+ $X2=3.235 $Y2=1.557
r44 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.235 $Y=1.765
+ $X2=3.235 $Y2=2.4
r45 1 11 24.7974 $w=3.11e-07 $l=2.75625e-07 $layer=POLY_cond $X=3.075 $Y=1.35
+ $X2=3.235 $Y2=1.557
r46 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.075 $Y=1.35
+ $X2=3.075 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_828_74# 1 2 7 9 12 14 16 18 19 21 24 25
+ 28 30 31 33 34 37 38 41 42 43 46 53 54 55 58 60 61 62 65 69
c199 65 0 1.41735e-19 $X=8.515 $Y=1.31
c200 61 0 8.50626e-20 $X=7.615 $Y=1.195
c201 53 0 2.22256e-19 $X=5.17 $Y=2.17
c202 33 0 1.21466e-19 $X=5.155 $Y=2.005
c203 12 0 1.1997e-19 $X=5.79 $Y=0.695
c204 7 0 1.03562e-19 $X=5.475 $Y=2.42
r205 69 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.515 $Y=1.39
+ $X2=8.515 $Y2=1.555
r206 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.515
+ $Y=1.39 $X2=8.515 $Y2=1.39
r207 65 68 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.515 $Y=1.31
+ $X2=8.515 $Y2=1.39
r208 61 76 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.615 $Y=1.195
+ $X2=7.48 $Y2=1.195
r209 60 63 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=7.65 $Y=1.195
+ $X2=7.65 $Y2=1.31
r210 60 62 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=1.195
+ $X2=7.65 $Y2=1.03
r211 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.615
+ $Y=1.195 $X2=7.615 $Y2=1.195
r212 58 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.84 $Y=1.21
+ $X2=5.84 $Y2=1.045
r213 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=1.21 $X2=5.84 $Y2=1.21
r214 55 57 16.8521 $w=2.57e-07 $l=3.55e-07 $layer=LI1_cond $X=5.915 $Y=0.855
+ $X2=5.915 $Y2=1.21
r215 53 72 51.947 $w=2.83e-07 $l=3.05e-07 $layer=POLY_cond $X=5.17 $Y=2.212
+ $X2=5.475 $Y2=2.212
r216 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.17
+ $Y=2.17 $X2=5.17 $Y2=2.17
r217 47 63 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.78 $Y=1.31
+ $X2=7.65 $Y2=1.31
r218 46 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.35 $Y=1.31
+ $X2=8.515 $Y2=1.31
r219 46 47 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.35 $Y=1.31
+ $X2=7.78 $Y2=1.31
r220 44 62 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.605 $Y=0.425
+ $X2=7.605 $Y2=1.03
r221 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.52 $Y=0.34
+ $X2=7.605 $Y2=0.425
r222 42 43 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.52 $Y=0.34
+ $X2=7.01 $Y2=0.34
r223 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.925 $Y=0.425
+ $X2=7.01 $Y2=0.34
r224 40 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.925 $Y=0.425
+ $X2=6.925 $Y2=0.77
r225 39 55 3.1561 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=0.855
+ $X2=5.915 $Y2=0.855
r226 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.84 $Y=0.855
+ $X2=6.925 $Y2=0.77
r227 38 39 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.84 $Y=0.855
+ $X2=6.08 $Y2=0.855
r228 37 55 5.43462 $w=2.57e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.995 $Y=0.77
+ $X2=5.915 $Y2=0.855
r229 36 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.995 $Y=0.425
+ $X2=5.995 $Y2=0.77
r230 35 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=0.34
+ $X2=5.155 $Y2=0.34
r231 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.91 $Y=0.34
+ $X2=5.995 $Y2=0.425
r232 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.91 $Y=0.34
+ $X2=5.24 $Y2=0.34
r233 33 52 0.582803 $w=3.14e-07 $l=1.5e-08 $layer=LI1_cond $X=5.155 $Y=2.072
+ $X2=5.17 $Y2=2.072
r234 33 49 18.0669 $w=3.14e-07 $l=4.65e-07 $layer=LI1_cond $X=5.155 $Y=2.072
+ $X2=4.69 $Y2=2.072
r235 32 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0.425
+ $X2=5.155 $Y2=0.34
r236 32 33 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=5.155 $Y=0.425
+ $X2=5.155 $Y2=2.005
r237 30 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=5.155 $Y2=0.34
r238 30 31 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=4.445 $Y2=0.34
r239 26 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.445 $Y2=0.34
r240 26 28 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.32 $Y2=0.515
r241 24 25 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.395 $Y=1.99
+ $X2=8.395 $Y2=2.14
r242 24 82 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.425 $Y=1.99
+ $X2=8.425 $Y2=1.555
r243 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.38 $Y=2.465
+ $X2=8.38 $Y2=2.75
r244 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.38 $Y=2.375
+ $X2=8.38 $Y2=2.465
r245 18 25 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=8.38 $Y=2.375
+ $X2=8.38 $Y2=2.14
r246 14 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.48 $Y=1.03
+ $X2=7.48 $Y2=1.195
r247 14 16 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.48 $Y=1.03
+ $X2=7.48 $Y2=0.645
r248 12 74 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.79 $Y=0.695
+ $X2=5.79 $Y2=1.045
r249 7 72 17.601 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.475 $Y=2.42
+ $X2=5.475 $Y2=2.212
r250 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.475 $Y=2.42
+ $X2=5.475 $Y2=2.705
r251 2 49 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=4.54
+ $Y=1.84 $X2=4.69 $Y2=2.01
r252 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_630_74# 1 2 9 11 13 15 16 20 22 25 26 28
+ 29 31 33 34 36 37 38 41 45 47 51 52 55 58 59 61 62 63 65 66 71 74 84
c202 71 0 5.59789e-20 $X=6.12 $Y=2.08
c203 61 0 2.69838e-19 $X=6.12 $Y=2.615
c204 58 0 6.34765e-20 $X=3.975 $Y=1.515
c205 41 0 3.61287e-20 $X=8.24 $Y=0.94
c206 38 0 1.21466e-19 $X=5.03 $Y=1.69
r207 75 84 18.4153 $w=3.01e-07 $l=1.15e-07 $layer=POLY_cond $X=7.73 $Y=1.822
+ $X2=7.845 $Y2=1.822
r208 74 77 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.73 $Y=1.765
+ $X2=7.73 $Y2=1.93
r209 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.73
+ $Y=1.765 $X2=7.73 $Y2=1.765
r210 68 71 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.965 $Y=2.08
+ $X2=6.12 $Y2=2.08
r211 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.965
+ $Y=2.08 $X2=5.965 $Y2=2.08
r212 65 77 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=7.65 $Y=2.615
+ $X2=7.65 $Y2=1.93
r213 62 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.565 $Y=2.7
+ $X2=7.65 $Y2=2.615
r214 62 63 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.565 $Y=2.7
+ $X2=6.205 $Y2=2.7
r215 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.12 $Y=2.615
+ $X2=6.205 $Y2=2.7
r216 60 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.12 $Y=2.245
+ $X2=6.12 $Y2=2.08
r217 60 61 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.12 $Y=2.245
+ $X2=6.12 $Y2=2.615
r218 59 80 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.975 $Y=1.515
+ $X2=3.975 $Y2=1.69
r219 59 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=1.515
+ $X2=3.975 $Y2=1.35
r220 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=1.515 $X2=3.975 $Y2=1.515
r221 56 58 20.888 $w=2.38e-07 $l=4.35e-07 $layer=LI1_cond $X=3.975 $Y=1.95
+ $X2=3.975 $Y2=1.515
r222 55 66 6.75802 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.975 $Y=1.47
+ $X2=3.975 $Y2=1.35
r223 55 58 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=3.975 $Y=1.47
+ $X2=3.975 $Y2=1.515
r224 53 66 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.94 $Y=1.18
+ $X2=3.94 $Y2=1.35
r225 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=1.095
+ $X2=3.94 $Y2=1.18
r226 51 52 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.855 $Y=1.095
+ $X2=3.455 $Y2=1.095
r227 47 56 6.82018 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=3.855 $Y=2.075
+ $X2=3.975 $Y2=1.95
r228 47 49 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=3.855 $Y=2.075
+ $X2=3.465 $Y2=2.075
r229 43 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.29 $Y=1.01
+ $X2=3.455 $Y2=1.095
r230 43 45 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.29 $Y=1.01
+ $X2=3.29 $Y2=0.515
r231 39 41 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=8.065 $Y=0.94
+ $X2=8.24 $Y2=0.94
r232 34 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.24 $Y=0.865
+ $X2=8.24 $Y2=0.94
r233 34 36 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.24 $Y=0.865
+ $X2=8.24 $Y2=0.58
r234 33 84 35.2292 $w=3.01e-07 $l=3.13247e-07 $layer=POLY_cond $X=8.065 $Y=1.6
+ $X2=7.845 $Y2=1.822
r235 32 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.065 $Y=1.015
+ $X2=8.065 $Y2=0.94
r236 32 33 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=8.065 $Y=1.015
+ $X2=8.065 $Y2=1.6
r237 29 84 19.0468 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.845 $Y=2.045
+ $X2=7.845 $Y2=1.822
r238 29 31 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.845 $Y=2.045
+ $X2=7.845 $Y2=2.54
r239 26 69 72.8652 $w=2.52e-07 $l=3.61801e-07 $layer=POLY_cond $X=6.01 $Y=2.42
+ $X2=5.965 $Y2=2.08
r240 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.01 $Y=2.42
+ $X2=6.01 $Y2=2.705
r241 25 69 2.81204 $w=3.3e-07 $l=8.75758e-08 $layer=POLY_cond $X=5.965 $Y=2.08
+ $X2=5.965 $Y2=2.08
r242 24 25 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=5.965 $Y=1.765
+ $X2=5.965 $Y2=2.08
r243 23 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.105 $Y=1.69
+ $X2=5.03 $Y2=1.69
r244 22 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.8 $Y=1.69
+ $X2=5.965 $Y2=1.765
r245 22 23 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.8 $Y=1.69
+ $X2=5.105 $Y2=1.69
r246 18 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.03 $Y=1.615
+ $X2=5.03 $Y2=1.69
r247 18 20 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=5.03 $Y=1.615
+ $X2=5.03 $Y2=0.695
r248 17 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.54 $Y=1.69
+ $X2=4.465 $Y2=1.69
r249 16 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.955 $Y=1.69
+ $X2=5.03 $Y2=1.69
r250 16 17 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.955 $Y=1.69
+ $X2=4.54 $Y2=1.69
r251 13 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.465 $Y=1.765
+ $X2=4.465 $Y2=1.69
r252 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.465 $Y=1.765
+ $X2=4.465 $Y2=2.4
r253 12 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.69
+ $X2=3.975 $Y2=1.69
r254 11 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.39 $Y=1.69
+ $X2=4.465 $Y2=1.69
r255 11 12 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.39 $Y=1.69
+ $X2=4.14 $Y2=1.69
r256 9 79 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.065 $Y=0.74
+ $X2=4.065 $Y2=1.35
r257 2 49 600 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=1.84 $X2=3.465 $Y2=2.115
r258 1 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.15
+ $Y=0.37 $X2=3.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_1243_48# 1 2 9 12 13 15 16 19 23 28 29 31
c70 12 0 5.59221e-20 $X=6.43 $Y=2.33
c71 9 0 1.1651e-19 $X=6.29 $Y=0.58
r72 28 29 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=7.252 $Y=2.28
+ $X2=7.252 $Y2=2.115
r73 25 31 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.265 $Y=1.405
+ $X2=7.265 $Y2=1.257
r74 25 29 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.265 $Y=1.405
+ $X2=7.265 $Y2=2.115
r75 21 31 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.265 $Y=1.11
+ $X2=7.265 $Y2=1.257
r76 21 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.265 $Y=1.11
+ $X2=7.265 $Y2=0.765
r77 19 34 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.397 $Y=1.24
+ $X2=6.397 $Y2=1.405
r78 19 33 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.397 $Y=1.24
+ $X2=6.397 $Y2=1.075
r79 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.415
+ $Y=1.24 $X2=6.415 $Y2=1.24
r80 16 31 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=1.257
+ $X2=7.265 $Y2=1.257
r81 16 18 29.8854 $w=2.93e-07 $l=7.65e-07 $layer=LI1_cond $X=7.18 $Y=1.257
+ $X2=6.415 $Y2=1.257
r82 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.43 $Y=2.42 $X2=6.43
+ $Y2=2.705
r83 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.43 $Y=2.33 $X2=6.43
+ $Y2=2.42
r84 12 34 359.556 $w=1.8e-07 $l=9.25e-07 $layer=POLY_cond $X=6.43 $Y=2.33
+ $X2=6.43 $Y2=1.405
r85 9 33 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.29 $Y=0.58
+ $X2=6.29 $Y2=1.075
r86 2 28 600 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_PDIFF $count=1 $X=7.125
+ $Y=2.12 $X2=7.29 $Y2=2.28
r87 1 23 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.37 $X2=7.265 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_1021_97# 1 2 9 11 13 15 18 21 24 26 27 29
c83 27 0 5.59221e-20 $X=5.685 $Y=2.475
c84 21 0 1.1651e-19 $X=5.575 $Y=0.695
r85 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.895
+ $Y=1.78 $X2=6.895 $Y2=1.78
r86 29 32 4.93904 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=6.87 $Y=1.66
+ $X2=6.87 $Y2=1.78
r87 26 27 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=5.685 $Y=2.705
+ $X2=5.685 $Y2=2.475
r88 21 23 8.98601 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.575 $Y=0.695
+ $X2=5.575 $Y2=0.875
r89 19 24 1.34256 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.675 $Y=1.66
+ $X2=5.542 $Y2=1.66
r90 18 29 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.73 $Y=1.66 $X2=6.87
+ $Y2=1.66
r91 18 19 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=6.73 $Y=1.66
+ $X2=5.675 $Y2=1.66
r92 16 24 5.16603 $w=1.7e-07 $l=1.06325e-07 $layer=LI1_cond $X=5.59 $Y=1.745
+ $X2=5.542 $Y2=1.66
r93 16 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.59 $Y=1.745
+ $X2=5.59 $Y2=2.475
r94 15 24 5.16603 $w=1.7e-07 $l=1.05924e-07 $layer=LI1_cond $X=5.495 $Y=1.575
+ $X2=5.542 $Y2=1.66
r95 15 23 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.495 $Y=1.575
+ $X2=5.495 $Y2=0.875
r96 11 33 52.3966 $w=3.56e-07 $l=3.17333e-07 $layer=POLY_cond $X=7.05 $Y=2.045
+ $X2=6.935 $Y2=1.78
r97 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.05 $Y=2.045
+ $X2=7.05 $Y2=2.54
r98 7 33 38.8573 $w=3.56e-07 $l=2.14942e-07 $layer=POLY_cond $X=7.05 $Y=1.615
+ $X2=6.935 $Y2=1.78
r99 7 9 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.05 $Y=1.615 $X2=7.05
+ $Y2=0.645
r100 2 26 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=5.55
+ $Y=2.495 $X2=5.7 $Y2=2.705
r101 1 21 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.485 $X2=5.575 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_1711_48# 1 2 7 9 10 11 12 14 16 17 19 21
+ 24 26 29 30 32 35 37 40 41 43 46 48 49 50 57 60 62 65 69 73 74
c164 11 0 1.41735e-19 $X=8.705 $Y=0.94
r165 69 71 11.5626 $w=3.88e-07 $l=2.65e-07 $layer=LI1_cond $X=9.755 $Y=0.62
+ $X2=9.755 $Y2=0.885
r166 63 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.95 $Y=1.465
+ $X2=9.865 $Y2=1.465
r167 63 65 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=9.95 $Y=1.465
+ $X2=10.445 $Y2=1.465
r168 62 73 6.11814 $w=2.6e-07 $l=2.61151e-07 $layer=LI1_cond $X=9.865 $Y=1.94
+ $X2=9.775 $Y2=2.16
r169 61 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.63
+ $X2=9.865 $Y2=1.465
r170 61 62 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.865 $Y=1.63
+ $X2=9.865 $Y2=1.94
r171 60 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.3
+ $X2=9.865 $Y2=1.465
r172 60 71 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.865 $Y=1.3
+ $X2=9.865 $Y2=0.885
r173 55 73 6.11814 $w=2.6e-07 $l=2.2e-07 $layer=LI1_cond $X=9.775 $Y=2.38
+ $X2=9.775 $Y2=2.16
r174 55 57 14.3232 $w=3.48e-07 $l=4.35e-07 $layer=LI1_cond $X=9.775 $Y=2.38
+ $X2=9.775 $Y2=2.815
r175 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.875
+ $Y=2.215 $X2=8.875 $Y2=2.215
r176 50 73 0.606672 $w=3.2e-07 $l=2.02793e-07 $layer=LI1_cond $X=9.6 $Y=2.22
+ $X2=9.775 $Y2=2.16
r177 50 52 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=9.6 $Y=2.22
+ $X2=8.875 $Y2=2.22
r178 44 49 18.8402 $w=1.65e-07 $l=8.35165e-08 $layer=POLY_cond $X=11.99 $Y=1.3
+ $X2=11.972 $Y2=1.375
r179 44 46 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=11.99 $Y=1.3
+ $X2=11.99 $Y2=0.81
r180 41 43 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.97 $Y=1.765
+ $X2=11.97 $Y2=2.34
r181 40 41 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.97 $Y=1.675
+ $X2=11.97 $Y2=1.765
r182 39 49 18.8402 $w=1.65e-07 $l=7.59934e-08 $layer=POLY_cond $X=11.97 $Y=1.45
+ $X2=11.972 $Y2=1.375
r183 39 40 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=11.97 $Y=1.45
+ $X2=11.97 $Y2=1.675
r184 38 48 13.2179 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=11.075 $Y=1.375
+ $X2=10.982 $Y2=1.375
r185 37 49 6.66866 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=11.88 $Y=1.375
+ $X2=11.972 $Y2=1.375
r186 37 38 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=11.88 $Y=1.375
+ $X2=11.075 $Y2=1.375
r187 33 48 10.9219 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=11 $Y=1.3
+ $X2=10.982 $Y2=1.375
r188 33 35 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11 $Y=1.3 $X2=11
+ $Y2=0.74
r189 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.98 $Y=1.765
+ $X2=10.98 $Y2=2.4
r190 29 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.98 $Y=1.675
+ $X2=10.98 $Y2=1.765
r191 28 48 10.9219 $w=1.8e-07 $l=7.59934e-08 $layer=POLY_cond $X=10.98 $Y=1.45
+ $X2=10.982 $Y2=1.375
r192 28 29 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=10.98 $Y=1.45
+ $X2=10.98 $Y2=1.675
r193 27 76 9.2281 $w=1.5e-07 $l=1.03e-07 $layer=POLY_cond $X=10.645 $Y=1.375
+ $X2=10.542 $Y2=1.375
r194 26 48 13.2179 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=10.89 $Y=1.375
+ $X2=10.982 $Y2=1.375
r195 26 27 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=10.89 $Y=1.375
+ $X2=10.645 $Y2=1.375
r196 22 76 21.2113 $w=1.97e-07 $l=8.7892e-08 $layer=POLY_cond $X=10.57 $Y=1.3
+ $X2=10.542 $Y2=1.375
r197 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.57 $Y=1.3
+ $X2=10.57 $Y2=0.74
r198 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=2.4
r199 17 19 76.2621 $w=1.97e-07 $l=3.05941e-07 $layer=POLY_cond $X=10.542
+ $Y=1.465 $X2=10.53 $Y2=1.765
r200 17 76 22.0203 $w=1.97e-07 $l=9e-08 $layer=POLY_cond $X=10.542 $Y=1.465
+ $X2=10.542 $Y2=1.375
r201 17 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.445
+ $Y=1.465 $X2=10.445 $Y2=1.465
r202 16 53 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=8.965 $Y=2.05
+ $X2=8.875 $Y2=2.215
r203 15 16 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=8.965 $Y=1.015
+ $X2=8.965 $Y2=2.05
r204 12 53 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=8.8 $Y=2.465
+ $X2=8.875 $Y2=2.215
r205 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.8 $Y=2.465 $X2=8.8
+ $Y2=2.75
r206 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.89 $Y=0.94
+ $X2=8.965 $Y2=1.015
r207 10 11 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=8.89 $Y=0.94
+ $X2=8.705 $Y2=0.94
r208 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.63 $Y=0.865
+ $X2=8.705 $Y2=0.94
r209 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.63 $Y=0.865 $X2=8.63
+ $Y2=0.58
r210 2 73 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.615
+ $Y=1.96 $X2=9.765 $Y2=2.105
r211 2 57 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=9.615
+ $Y=1.96 $X2=9.765 $Y2=2.815
r212 1 69 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=9.585
+ $Y=0.37 $X2=9.725 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_1511_74# 1 2 9 11 12 14 17 19 23 25 26 28
+ 29 32 34 35 38 42 45
c110 35 0 3.61287e-20 $X=8.935 $Y=0.97
c111 32 0 8.50626e-20 $X=8.025 $Y=0.58
r112 42 46 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.455 $Y=1.385
+ $X2=9.455 $Y2=1.55
r113 42 45 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.455 $Y=1.385
+ $X2=9.455 $Y2=1.22
r114 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.445
+ $Y=1.385 $X2=9.445 $Y2=1.385
r115 38 41 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=9.445 $Y=1.14
+ $X2=9.445 $Y2=1.385
r116 35 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.935 $Y=0.97
+ $X2=8.935 $Y2=1.14
r117 32 33 17.365 $w=2.74e-07 $l=3.9e-07 $layer=LI1_cond $X=8.025 $Y=0.58
+ $X2=8.025 $Y2=0.97
r118 30 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.02 $Y=1.14
+ $X2=8.935 $Y2=1.14
r119 29 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.28 $Y=1.14
+ $X2=9.445 $Y2=1.14
r120 29 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.28 $Y=1.14
+ $X2=9.02 $Y2=1.14
r121 27 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=1.225
+ $X2=8.935 $Y2=1.14
r122 27 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.935 $Y=1.225
+ $X2=8.935 $Y2=1.72
r123 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.85 $Y=1.805
+ $X2=8.935 $Y2=1.72
r124 25 26 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=8.85 $Y=1.805
+ $X2=8.235 $Y2=1.805
r125 24 33 3.52985 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=0.97
+ $X2=8.025 $Y2=0.97
r126 23 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=0.97
+ $X2=8.935 $Y2=0.97
r127 23 24 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.85 $Y=0.97
+ $X2=8.19 $Y2=0.97
r128 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.15 $Y=1.89
+ $X2=8.235 $Y2=1.805
r129 21 34 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.15 $Y=1.89
+ $X2=8.15 $Y2=2.1
r130 17 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=2.265
+ $X2=8.07 $Y2=2.1
r131 17 19 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=8.07 $Y=2.265
+ $X2=8.07 $Y2=2.815
r132 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.54 $Y=1.885
+ $X2=9.54 $Y2=2.46
r133 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.54 $Y=1.795
+ $X2=9.54 $Y2=1.885
r134 11 46 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=9.54 $Y=1.795
+ $X2=9.54 $Y2=1.55
r135 9 45 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.51 $Y=0.74 $X2=9.51
+ $Y2=1.22
r136 2 19 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=7.92
+ $Y=2.12 $X2=8.07 $Y2=2.815
r137 2 17 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.92
+ $Y=2.12 $X2=8.07 $Y2=2.265
r138 1 32 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=7.555
+ $Y=0.37 $X2=8.025 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_2322_368# 1 2 7 9 12 16 18 20 23 27 33 36
+ 40
c73 27 0 1.47924e-19 $X=11.745 $Y=1.985
r74 37 38 0.610127 $w=3.95e-07 $l=5e-09 $layer=POLY_cond $X=12.495 $Y=1.542
+ $X2=12.5 $Y2=1.542
r75 34 40 45.7595 $w=3.95e-07 $l=3.75e-07 $layer=POLY_cond $X=12.57 $Y=1.542
+ $X2=12.945 $Y2=1.542
r76 34 38 8.54177 $w=3.95e-07 $l=7e-08 $layer=POLY_cond $X=12.57 $Y=1.542
+ $X2=12.5 $Y2=1.542
r77 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.57
+ $Y=1.485 $X2=12.57 $Y2=1.485
r78 31 36 1.50311 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=11.94 $Y=1.485
+ $X2=11.76 $Y2=1.485
r79 31 33 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=11.94 $Y=1.485
+ $X2=12.57 $Y2=1.485
r80 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=11.745 $Y=1.985
+ $X2=11.745 $Y2=2.695
r81 25 36 4.97762 $w=3.45e-07 $l=1.72337e-07 $layer=LI1_cond $X=11.745 $Y=1.65
+ $X2=11.76 $Y2=1.485
r82 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.745 $Y=1.65
+ $X2=11.745 $Y2=1.985
r83 21 36 4.97762 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=11.76 $Y=1.32
+ $X2=11.76 $Y2=1.485
r84 21 23 20.9681 $w=3.58e-07 $l=6.55e-07 $layer=LI1_cond $X=11.76 $Y=1.32
+ $X2=11.76 $Y2=0.665
r85 18 40 25.5547 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=12.945 $Y=1.765
+ $X2=12.945 $Y2=1.542
r86 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.945 $Y=1.765
+ $X2=12.945 $Y2=2.4
r87 14 40 25.5547 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=12.945 $Y=1.32
+ $X2=12.945 $Y2=1.542
r88 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.945 $Y=1.32
+ $X2=12.945 $Y2=0.76
r89 10 38 25.5547 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=12.5 $Y=1.32
+ $X2=12.5 $Y2=1.542
r90 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.5 $Y=1.32
+ $X2=12.5 $Y2=0.76
r91 7 37 25.5547 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=12.495 $Y=1.765
+ $X2=12.495 $Y2=1.542
r92 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.495 $Y=1.765
+ $X2=12.495 $Y2=2.4
r93 2 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=11.61
+ $Y=1.84 $X2=11.745 $Y2=2.695
r94 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.61
+ $Y=1.84 $X2=11.745 $Y2=1.985
r95 1 23 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=11.63
+ $Y=0.49 $X2=11.775 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 53
+ 56 60 64 66 69 70 72 73 75 78 82 83 85 97 108 116 120 125 131 134 137 140 144
c166 30 0 1.92539e-19 $X=0.89 $Y=2.41
r167 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r168 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r169 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r170 134 135 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r171 131 132 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r172 129 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r173 129 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r174 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r175 126 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.355 $Y=3.33
+ $X2=12.23 $Y2=3.33
r176 126 128 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.355 $Y=3.33
+ $X2=12.72 $Y2=3.33
r177 125 143 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=13.222 $Y2=3.33
r178 125 128 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=12.72 $Y2=3.33
r179 124 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r180 124 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r181 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r182 121 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.205 $Y2=3.33
r183 121 123 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.76 $Y2=3.33
r184 120 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.105 $Y=3.33
+ $X2=12.23 $Y2=3.33
r185 120 123 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.105 $Y=3.33
+ $X2=11.76 $Y2=3.33
r186 119 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r187 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r188 116 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=11.205 $Y2=3.33
r189 116 118 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=10.8 $Y2=3.33
r190 115 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r191 115 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r192 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r193 112 134 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.145 $Y2=3.33
r194 112 114 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.84 $Y2=3.33
r195 111 135 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r196 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r197 108 134 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=9.145 $Y2=3.33
r198 108 110 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=6.96 $Y2=3.33
r199 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r200 104 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r201 104 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r202 103 106 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r203 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r204 101 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.24 $Y2=3.33
r205 101 103 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.56 $Y2=3.33
r206 100 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r207 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r208 97 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=4.24 $Y2=3.33
r209 97 99 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=3.12 $Y2=3.33
r210 96 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r211 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r212 93 96 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r213 92 95 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r214 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r215 89 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r216 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r217 85 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r218 85 107 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r219 82 114 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=9.84 $Y2=3.33
r220 82 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=10.265 $Y2=3.33
r221 81 118 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=10.39 $Y=3.33
+ $X2=10.8 $Y2=3.33
r222 81 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.39 $Y=3.33
+ $X2=10.265 $Y2=3.33
r223 79 110 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.905 $Y=3.33
+ $X2=6.96 $Y2=3.33
r224 78 106 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.575 $Y=3.33
+ $X2=6.48 $Y2=3.33
r225 77 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=3.33
+ $X2=6.905 $Y2=3.33
r226 77 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=3.33
+ $X2=6.575 $Y2=3.33
r227 75 77 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=6.74 $Y=3.04
+ $X2=6.74 $Y2=3.33
r228 72 95 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=3.33 $X2=2.64
+ $Y2=3.33
r229 72 73 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.88 $Y2=3.33
r230 71 99 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.09 $Y=3.33 $X2=3.12
+ $Y2=3.33
r231 71 73 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.09 $Y=3.33
+ $X2=2.88 $Y2=3.33
r232 69 88 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r233 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r234 68 92 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r235 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r236 64 143 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.222 $Y2=3.33
r237 64 66 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=2.405
r238 60 63 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.23 $Y=1.985
+ $X2=12.23 $Y2=2.815
r239 58 140 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.23 $Y=3.245
+ $X2=12.23 $Y2=3.33
r240 58 63 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.23 $Y=3.245
+ $X2=12.23 $Y2=2.815
r241 56 84 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=11.245 $Y=1.985
+ $X2=11.245 $Y2=2.14
r242 51 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.205 $Y=3.245
+ $X2=11.205 $Y2=3.33
r243 51 53 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=11.205 $Y=3.245
+ $X2=11.205 $Y2=2.4
r244 50 84 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.205 $Y=2.305
+ $X2=11.205 $Y2=2.14
r245 50 53 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=11.205 $Y=2.305
+ $X2=11.205 $Y2=2.4
r246 46 49 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.265 $Y=1.985
+ $X2=10.265 $Y2=2.815
r247 44 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=3.245
+ $X2=10.265 $Y2=3.33
r248 44 49 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.265 $Y=3.245
+ $X2=10.265 $Y2=2.815
r249 40 134 2.39972 $w=5.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=3.33
r250 40 42 9.02305 $w=5.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=2.815
r251 36 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=3.245
+ $X2=4.24 $Y2=3.33
r252 36 38 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.24 $Y=3.245
+ $X2=4.24 $Y2=2.805
r253 32 73 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=3.33
r254 32 34 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=2.875
r255 28 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=3.33
r256 28 30 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=2.41
r257 9 66 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=13.02
+ $Y=1.84 $X2=13.17 $Y2=2.405
r258 8 63 600 $w=1.7e-07 $l=1.08167e-06 $layer=licon1_PDIFF $count=1 $X=12.045
+ $Y=1.84 $X2=12.27 $Y2=2.815
r259 8 60 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=12.045
+ $Y=1.84 $X2=12.27 $Y2=1.985
r260 7 56 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.055
+ $Y=1.84 $X2=11.205 $Y2=1.985
r261 7 53 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=11.055
+ $Y=1.84 $X2=11.205 $Y2=2.4
r262 6 49 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.305 $Y2=2.815
r263 6 46 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.305 $Y2=1.985
r264 5 42 600 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_PDIFF $count=1 $X=8.875
+ $Y=2.54 $X2=9.145 $Y2=2.815
r265 4 75 600 $w=1.7e-07 $l=6.51997e-07 $layer=licon1_PDIFF $count=1 $X=6.505
+ $Y=2.495 $X2=6.74 $Y2=3.04
r266 3 38 600 $w=1.7e-07 $l=1.03496e-06 $layer=licon1_PDIFF $count=1 $X=4.095
+ $Y=1.84 $X2=4.24 $Y2=2.805
r267 2 34 600 $w=1.7e-07 $l=7.36818e-07 $layer=licon1_PDIFF $count=1 $X=2.6
+ $Y=2.265 $X2=2.88 $Y2=2.875
r268 1 30 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.74
+ $Y=2.265 $X2=0.89 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%A_301_74# 1 2 3 4 13 19 22 23 24 26 27 30
+ 31 32 35 37 38 40 41 43
c122 24 0 6.78066e-20 $X=2.415 $Y=1.435
r123 43 46 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=5.21 $Y=2.58
+ $X2=5.21 $Y2=2.715
r124 38 42 23.0691 $w=2.14e-07 $l=4.25335e-07 $layer=LI1_cond $X=4.745 $Y=2.58
+ $X2=4.35 $Y2=2.517
r125 37 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.085 $Y=2.58
+ $X2=5.21 $Y2=2.58
r126 37 38 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.085 $Y=2.58
+ $X2=4.745 $Y2=2.58
r127 33 35 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=4.775 $Y=1.48
+ $X2=4.775 $Y2=0.76
r128 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.65 $Y=1.565
+ $X2=4.775 $Y2=1.48
r129 31 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.65 $Y=1.565
+ $X2=4.435 $Y2=1.565
r130 30 42 2.08775 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=4.35 $Y=2.37
+ $X2=4.35 $Y2=2.517
r131 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=1.65
+ $X2=4.435 $Y2=1.565
r132 29 30 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.35 $Y=1.65
+ $X2=4.35 $Y2=2.37
r133 28 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=2.455
+ $X2=3.01 $Y2=2.455
r134 27 42 5.39616 $w=2.14e-07 $l=1.11781e-07 $layer=LI1_cond $X=4.265 $Y=2.455
+ $X2=4.35 $Y2=2.517
r135 27 28 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.265 $Y=2.455
+ $X2=3.095 $Y2=2.455
r136 26 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=2.37
+ $X2=3.01 $Y2=2.455
r137 25 26 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=3.01 $Y=1.52
+ $X2=3.01 $Y2=2.37
r138 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.925 $Y=1.435
+ $X2=3.01 $Y2=1.52
r139 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.925 $Y=1.435
+ $X2=2.415 $Y2=1.435
r140 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.33 $Y=1.35
+ $X2=2.415 $Y2=1.435
r141 21 22 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.33 $Y=0.64
+ $X2=2.33 $Y2=1.35
r142 20 40 4.88517 $w=1.7e-07 $l=1.79374e-07 $layer=LI1_cond $X=1.98 $Y=2.455
+ $X2=1.815 $Y2=2.425
r143 19 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=2.455
+ $X2=3.01 $Y2=2.455
r144 19 20 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=2.925 $Y=2.455
+ $X2=1.98 $Y2=2.455
r145 13 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.245 $Y=0.515
+ $X2=2.33 $Y2=0.64
r146 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.245 $Y=0.515
+ $X2=1.8 $Y2=0.515
r147 4 46 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=5.105
+ $Y=2.495 $X2=5.25 $Y2=2.715
r148 3 40 300 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=2 $X=1.61
+ $Y=2.265 $X2=1.815 $Y2=2.41
r149 2 35 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=4.68
+ $Y=0.485 $X2=4.815 $Y2=0.76
r150 1 15 182 $w=1.7e-07 $l=3.76298e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.37 $X2=1.8 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%Q 1 2 9 15 16 17 18 29
r39 22 29 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=10.785 $Y=0.965
+ $X2=10.785 $Y2=0.925
r40 18 31 7.69388 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=10.785 $Y=0.987
+ $X2=10.785 $Y2=1.13
r41 18 22 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=10.785 $Y=0.987
+ $X2=10.785 $Y2=0.965
r42 18 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=10.785 $Y=0.902
+ $X2=10.785 $Y2=0.925
r43 17 18 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=10.785 $Y=0.515
+ $X2=10.785 $Y2=0.902
r44 15 16 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=10.77 $Y=1.8
+ $X2=10.77 $Y2=1.97
r45 15 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.865 $Y=1.8
+ $X2=10.865 $Y2=1.13
r46 9 11 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.715 $Y=1.985
+ $X2=10.715 $Y2=2.815
r47 9 16 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=10.715 $Y=1.985
+ $X2=10.715 $Y2=1.97
r48 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.755 $Y2=2.815
r49 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.755 $Y2=1.985
r50 1 17 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.645
+ $Y=0.37 $X2=10.785 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%Q_N 1 2 7 13 16 17 18
r29 30 31 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=13.195 $Y2=1.985
r30 27 30 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=12.695 $Y=1.985
+ $X2=12.72 $Y2=1.985
r31 22 31 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.82
+ $X2=13.195 $Y2=1.985
r32 18 31 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=13.2 $Y=1.985
+ $X2=13.195 $Y2=1.985
r33 17 22 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=13.195 $Y=1.665
+ $X2=13.195 $Y2=1.82
r34 16 17 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=13.195 $Y=1.295
+ $X2=13.195 $Y2=1.665
r35 15 16 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=13.195 $Y=1.15
+ $X2=13.195 $Y2=1.295
r36 11 27 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.695 $Y=2.15
+ $X2=12.695 $Y2=1.985
r37 11 13 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=12.695 $Y=2.15
+ $X2=12.695 $Y2=2.4
r38 7 15 6.82018 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=13.075 $Y=1.025
+ $X2=13.195 $Y2=1.15
r39 7 9 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=13.075 $Y=1.025
+ $X2=12.72 $Y2=1.025
r40 2 30 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.57
+ $Y=1.84 $X2=12.72 $Y2=1.985
r41 2 13 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=12.57
+ $Y=1.84 $X2=12.72 $Y2=2.4
r42 1 9 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=12.575
+ $Y=0.39 $X2=12.72 $Y2=0.985
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_2%VGND 1 2 3 4 5 6 7 8 9 32 36 42 46 50 54 59
+ 62 64 66 69 70 72 73 74 75 87 94 102 107 112 117 123 126 130 136 139 142 146
c159 46 0 1.1997e-19 $X=6.505 $Y=0.515
r160 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r161 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r162 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r163 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r164 130 133 9.0127 $w=7.08e-07 $l=5.35e-07 $layer=LI1_cond $X=9.035 $Y=0
+ $X2=9.035 $Y2=0.535
r165 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r166 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r167 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r168 121 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r169 121 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r170 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r171 118 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.45 $Y=0
+ $X2=12.285 $Y2=0
r172 118 120 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12.45 $Y=0
+ $X2=12.72 $Y2=0
r173 117 145 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.995 $Y=0
+ $X2=13.217 $Y2=0
r174 117 120 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.995 $Y=0
+ $X2=12.72 $Y2=0
r175 116 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r176 116 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r177 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r178 113 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.38 $Y=0
+ $X2=11.255 $Y2=0
r179 113 115 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.38 $Y=0
+ $X2=11.76 $Y2=0
r180 112 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.12 $Y=0
+ $X2=12.285 $Y2=0
r181 112 115 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=12.12 $Y=0
+ $X2=11.76 $Y2=0
r182 111 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r183 111 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r184 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r185 108 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=0
+ $X2=10.285 $Y2=0
r186 108 110 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=10.45 $Y=0
+ $X2=10.8 $Y2=0
r187 107 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.13 $Y=0
+ $X2=11.255 $Y2=0
r188 107 110 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=11.13 $Y=0
+ $X2=10.8 $Y2=0
r189 106 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r190 106 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r191 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r192 103 130 9.41505 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=9.39 $Y=0
+ $X2=9.035 $Y2=0
r193 103 105 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.39 $Y=0
+ $X2=9.84 $Y2=0
r194 102 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.12 $Y=0
+ $X2=10.285 $Y2=0
r195 102 105 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.12 $Y=0
+ $X2=9.84 $Y2=0
r196 101 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r197 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r198 98 101 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.4 $Y2=0
r199 97 100 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r200 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r201 95 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=6.505 $Y2=0
r202 95 97 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.96
+ $Y2=0
r203 94 130 9.41505 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=8.68 $Y=0
+ $X2=9.035 $Y2=0
r204 94 100 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.68 $Y=0 $X2=8.4
+ $Y2=0
r205 93 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r206 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r207 90 93 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r208 89 92 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r209 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r210 87 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=0
+ $X2=6.505 $Y2=0
r211 87 92 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.34 $Y=0 $X2=6
+ $Y2=0
r212 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r213 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r214 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r215 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r216 80 83 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r217 80 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r218 79 82 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r219 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r220 77 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0
+ $X2=0.825 $Y2=0
r221 77 79 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r222 75 98 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.96 $Y2=0
r223 75 127 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.48 $Y2=0
r224 72 85 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r225 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.85
+ $Y2=0
r226 71 89 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.08
+ $Y2=0
r227 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.85
+ $Y2=0
r228 69 82 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.64
+ $Y2=0
r229 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.82
+ $Y2=0
r230 68 85 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.6
+ $Y2=0
r231 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.82
+ $Y2=0
r232 64 145 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=13.16 $Y=0.085
+ $X2=13.217 $Y2=0
r233 64 66 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=13.16 $Y=0.085
+ $X2=13.16 $Y2=0.55
r234 62 74 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=12.25 $Y=0.985
+ $X2=12.25 $Y2=0.73
r235 57 74 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.285 $Y=0.565
+ $X2=12.285 $Y2=0.73
r236 57 59 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=12.285 $Y=0.565
+ $X2=12.285 $Y2=0.55
r237 56 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.285 $Y=0.085
+ $X2=12.285 $Y2=0
r238 56 59 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=12.285 $Y=0.085
+ $X2=12.285 $Y2=0.55
r239 52 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.255 $Y=0.085
+ $X2=11.255 $Y2=0
r240 52 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.255 $Y=0.085
+ $X2=11.255 $Y2=0.515
r241 48 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0
r242 48 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.515
r243 44 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0.085
+ $X2=6.505 $Y2=0
r244 44 46 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.505 $Y=0.085
+ $X2=6.505 $Y2=0.515
r245 40 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0
r246 40 42 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0.595
r247 36 38 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.82 $Y=0.515
+ $X2=2.82 $Y2=0.965
r248 34 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=0.085
+ $X2=2.82 $Y2=0
r249 34 36 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.82 $Y=0.085
+ $X2=2.82 $Y2=0.515
r250 30 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r251 30 32 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.54
r252 9 66 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=13.02
+ $Y=0.39 $X2=13.16 $Y2=0.55
r253 8 62 182 $w=1.7e-07 $l=5.82301e-07 $layer=licon1_NDIFF $count=1 $X=12.065
+ $Y=0.49 $X2=12.255 $Y2=0.985
r254 8 59 182 $w=1.7e-07 $l=2.48193e-07 $layer=licon1_NDIFF $count=1 $X=12.065
+ $Y=0.49 $X2=12.285 $Y2=0.55
r255 7 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.075
+ $Y=0.37 $X2=11.215 $Y2=0.515
r256 6 50 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.14
+ $Y=0.37 $X2=10.285 $Y2=0.515
r257 5 133 91 $w=1.7e-07 $l=6.6742e-07 $layer=licon1_NDIFF $count=2 $X=8.705
+ $Y=0.37 $X2=9.295 $Y2=0.535
r258 4 46 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.365
+ $Y=0.37 $X2=6.505 $Y2=0.515
r259 3 42 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.37 $X2=3.85 $Y2=0.595
r260 2 38 182 $w=1.7e-07 $l=6.96366e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.37 $X2=2.86 $Y2=0.965
r261 2 36 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.37 $X2=2.86 $Y2=0.515
r262 1 32 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.37 $X2=0.825 $Y2=0.54
.ends

