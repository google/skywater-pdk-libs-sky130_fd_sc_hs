# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__o2bb2a_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__o2bb2a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.475000 2.865000 1.805000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.475000 2.325000 1.805000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.570000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.810000 1.450000 1.285000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425000 1.820000 3.770000 2.980000 ;
        RECT 3.430000 0.350000 3.770000 1.130000 ;
        RECT 3.600000 1.130000 3.770000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.110000 ;
      RECT 0.115000  1.110000 1.305000 1.280000 ;
      RECT 0.120000  1.950000 0.450000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.940000 ;
      RECT 1.050000  1.950000 1.380000 2.395000 ;
      RECT 1.050000  2.395000 3.255000 2.565000 ;
      RECT 1.050000  2.565000 1.380000 2.980000 ;
      RECT 1.055000  0.350000 1.305000 1.110000 ;
      RECT 1.455000  1.450000 1.785000 1.780000 ;
      RECT 1.475000  0.255000 2.715000 0.425000 ;
      RECT 1.475000  0.425000 1.805000 0.965000 ;
      RECT 1.585000  2.735000 1.940000 3.245000 ;
      RECT 1.615000  1.135000 2.375000 1.305000 ;
      RECT 1.615000  1.305000 1.785000 1.450000 ;
      RECT 1.615000  1.780000 1.785000 1.975000 ;
      RECT 1.615000  1.975000 2.565000 2.225000 ;
      RECT 2.045000  0.595000 2.375000 1.135000 ;
      RECT 2.545000  0.425000 2.715000 1.135000 ;
      RECT 2.545000  1.135000 3.255000 1.305000 ;
      RECT 2.770000  2.735000 3.220000 3.245000 ;
      RECT 2.885000  0.085000 3.215000 0.965000 ;
      RECT 3.085000  1.305000 3.430000 1.635000 ;
      RECT 3.085000  1.635000 3.255000 2.395000 ;
      RECT 3.940000  0.085000 4.190000 1.130000 ;
      RECT 3.955000  1.820000 4.205000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o2bb2a_2
