* File: sky130_fd_sc_hs__a222oi_2.pxi.spice
* Created: Tue Sep  1 19:51:00 2020
* 
x_PM_SKY130_FD_SC_HS__A222OI_2%C2 N_C2_c_126_n N_C2_c_136_n N_C2_M1009_g
+ N_C2_M1014_g N_C2_c_137_n N_C2_M1012_g N_C2_M1016_g N_C2_c_128_n N_C2_c_129_n
+ N_C2_c_130_n N_C2_c_139_n N_C2_c_140_n N_C2_c_131_n N_C2_c_132_n C2
+ N_C2_c_134_n PM_SKY130_FD_SC_HS__A222OI_2%C2
x_PM_SKY130_FD_SC_HS__A222OI_2%C1 N_C1_c_225_n N_C1_M1007_g N_C1_M1002_g
+ N_C1_c_220_n N_C1_c_221_n N_C1_c_228_n N_C1_M1010_g N_C1_M1017_g N_C1_c_229_n
+ C1 N_C1_c_224_n PM_SKY130_FD_SC_HS__A222OI_2%C1
x_PM_SKY130_FD_SC_HS__A222OI_2%B1 N_B1_M1022_g N_B1_c_282_n N_B1_M1005_g
+ N_B1_c_283_n N_B1_M1019_g N_B1_M1023_g N_B1_c_285_n N_B1_c_291_n N_B1_c_292_n
+ N_B1_c_331_p N_B1_c_293_n N_B1_c_286_n B1 N_B1_c_287_n
+ PM_SKY130_FD_SC_HS__A222OI_2%B1
x_PM_SKY130_FD_SC_HS__A222OI_2%B2 N_B2_M1015_g N_B2_c_376_n N_B2_c_382_n
+ N_B2_M1020_g N_B2_c_377_n N_B2_c_384_n N_B2_M1021_g N_B2_c_378_n N_B2_M1018_g
+ B2 N_B2_c_379_n N_B2_c_380_n PM_SKY130_FD_SC_HS__A222OI_2%B2
x_PM_SKY130_FD_SC_HS__A222OI_2%A1 N_A1_M1011_g N_A1_c_442_n N_A1_M1006_g
+ N_A1_M1013_g N_A1_c_444_n N_A1_M1008_g N_A1_c_449_n N_A1_c_450_n N_A1_c_494_p
+ N_A1_c_451_n N_A1_c_445_n A1 N_A1_c_446_n PM_SKY130_FD_SC_HS__A222OI_2%A1
x_PM_SKY130_FD_SC_HS__A222OI_2%A2 N_A2_c_532_n N_A2_M1003_g N_A2_M1000_g
+ N_A2_c_533_n N_A2_M1004_g N_A2_M1001_g A2 N_A2_c_531_n
+ PM_SKY130_FD_SC_HS__A222OI_2%A2
x_PM_SKY130_FD_SC_HS__A222OI_2%Y N_Y_M1002_s N_Y_M1022_s N_Y_M1023_s N_Y_M1013_s
+ N_Y_M1009_s N_Y_M1007_s N_Y_M1012_s N_Y_c_584_n N_Y_c_585_n N_Y_c_604_n
+ N_Y_c_685_p N_Y_c_609_n N_Y_c_586_n N_Y_c_587_n N_Y_c_588_n N_Y_c_589_n
+ N_Y_c_590_n N_Y_c_591_n N_Y_c_592_n N_Y_c_619_n N_Y_c_620_n N_Y_c_622_n
+ N_Y_c_595_n Y Y Y PM_SKY130_FD_SC_HS__A222OI_2%Y
x_PM_SKY130_FD_SC_HS__A222OI_2%A_116_392# N_A_116_392#_M1009_d
+ N_A_116_392#_M1010_d N_A_116_392#_M1005_s N_A_116_392#_M1021_s
+ N_A_116_392#_c_738_n N_A_116_392#_c_732_n N_A_116_392#_c_733_n
+ N_A_116_392#_c_740_n N_A_116_392#_c_734_n N_A_116_392#_c_735_n
+ N_A_116_392#_c_736_n N_A_116_392#_c_737_n
+ PM_SKY130_FD_SC_HS__A222OI_2%A_116_392#
x_PM_SKY130_FD_SC_HS__A222OI_2%A_515_392# N_A_515_392#_M1005_d
+ N_A_515_392#_M1020_d N_A_515_392#_M1019_d N_A_515_392#_M1003_d
+ N_A_515_392#_M1008_d N_A_515_392#_c_796_n N_A_515_392#_c_839_n
+ N_A_515_392#_c_800_n N_A_515_392#_c_791_n N_A_515_392#_c_817_n
+ N_A_515_392#_c_792_n N_A_515_392#_c_821_n N_A_515_392#_c_793_n
+ N_A_515_392#_c_842_n N_A_515_392#_c_794_n N_A_515_392#_c_828_n
+ N_A_515_392#_c_795_n PM_SKY130_FD_SC_HS__A222OI_2%A_515_392#
x_PM_SKY130_FD_SC_HS__A222OI_2%VPWR N_VPWR_M1006_s N_VPWR_M1004_s N_VPWR_c_870_n
+ N_VPWR_c_871_n VPWR N_VPWR_c_872_n N_VPWR_c_873_n N_VPWR_c_874_n
+ N_VPWR_c_869_n N_VPWR_c_876_n N_VPWR_c_877_n PM_SKY130_FD_SC_HS__A222OI_2%VPWR
x_PM_SKY130_FD_SC_HS__A222OI_2%VGND N_VGND_M1014_d N_VGND_M1016_d N_VGND_M1015_d
+ N_VGND_M1000_d N_VGND_c_940_n N_VGND_c_941_n N_VGND_c_942_n N_VGND_c_943_n
+ VGND N_VGND_c_944_n N_VGND_c_945_n N_VGND_c_946_n N_VGND_c_947_n
+ N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n
+ PM_SKY130_FD_SC_HS__A222OI_2%VGND
x_PM_SKY130_FD_SC_HS__A222OI_2%A_137_74# N_A_137_74#_M1014_s N_A_137_74#_M1017_d
+ N_A_137_74#_c_1029_n PM_SKY130_FD_SC_HS__A222OI_2%A_137_74#
x_PM_SKY130_FD_SC_HS__A222OI_2%A_593_74# N_A_593_74#_M1022_d N_A_593_74#_M1018_s
+ N_A_593_74#_c_1044_n N_A_593_74#_c_1042_n N_A_593_74#_c_1043_n
+ PM_SKY130_FD_SC_HS__A222OI_2%A_593_74#
x_PM_SKY130_FD_SC_HS__A222OI_2%A_981_74# N_A_981_74#_M1011_d N_A_981_74#_M1001_s
+ N_A_981_74#_c_1068_n N_A_981_74#_c_1075_n N_A_981_74#_c_1071_n
+ N_A_981_74#_c_1072_n N_A_981_74#_c_1069_n
+ PM_SKY130_FD_SC_HS__A222OI_2%A_981_74#
cc_1 VNB N_C2_c_126_n 0.0104319f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.795
cc_2 VNB N_C2_M1014_g 0.0214368f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_3 VNB N_C2_c_128_n 0.0207721f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.13
cc_4 VNB N_C2_c_129_n 0.0298256f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.635
cc_5 VNB N_C2_c_130_n 0.00280946f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_6 VNB N_C2_c_131_n 0.00263864f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_7 VNB N_C2_c_132_n 0.0188881f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_8 VNB C2 0.00453826f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_9 VNB N_C2_c_134_n 0.0330468f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.33
cc_10 VNB N_C1_M1002_g 0.0197442f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_11 VNB N_C1_c_220_n 0.00871426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C1_c_221_n 0.00871368f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=2.46
cc_13 VNB N_C1_M1017_g 0.0196961f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.13
cc_14 VNB C1 0.00139126f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.665
cc_15 VNB N_C1_c_224_n 0.0367937f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.33
cc_16 VNB N_B1_M1022_g 0.0415299f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_17 VNB N_B1_c_282_n 0.0188732f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_18 VNB N_B1_c_283_n 0.0166227f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_19 VNB N_B1_M1023_g 0.0345024f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=1.13
cc_20 VNB N_B1_c_285_n 0.00340496f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_21 VNB N_B1_c_286_n 0.00354957f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_22 VNB N_B1_c_287_n 0.00188639f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.165
cc_23 VNB N_B2_M1015_g 0.0261081f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_24 VNB N_B2_c_376_n 0.00348647f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_25 VNB N_B2_c_377_n 0.00359827f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=2.46
cc_26 VNB N_B2_c_378_n 0.0165083f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_27 VNB N_B2_c_379_n 0.00359946f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_28 VNB N_B2_c_380_n 0.0730061f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_29 VNB N_A1_M1011_g 0.0352532f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_30 VNB N_A1_c_442_n 0.0159606f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_31 VNB N_A1_M1013_g 0.0442873f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=1.885
cc_32 VNB N_A1_c_444_n 0.0204176f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=2.46
cc_33 VNB N_A1_c_445_n 0.00360097f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_34 VNB N_A1_c_446_n 0.0124003f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.33
cc_35 VNB N_A2_M1000_g 0.0342909f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_36 VNB N_A2_M1001_g 0.0328015f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=1.13
cc_37 VNB A2 0.00102026f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_38 VNB N_A2_c_531_n 0.0257392f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.75
cc_39 VNB N_Y_c_584_n 0.0315443f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.665
cc_40 VNB N_Y_c_585_n 0.00803133f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_41 VNB N_Y_c_586_n 0.00739598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_587_n 0.0077195f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.495
cc_43 VNB N_Y_c_588_n 0.0166262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_589_n 0.0234737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_590_n 0.0021982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_591_n 0.0321153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_592_n 0.0318202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VPWR_c_869_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.33
cc_49 VNB N_VGND_c_940_n 0.01289f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=1.13
cc_50 VNB N_VGND_c_941_n 0.0246219f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_51 VNB N_VGND_c_942_n 0.0128186f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.495
cc_52 VNB N_VGND_c_943_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.665
cc_53 VNB N_VGND_c_944_n 0.0378216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_945_n 0.0317955f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.495
cc_55 VNB N_VGND_c_946_n 0.0415162f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.495
cc_56 VNB N_VGND_c_947_n 0.0299361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_948_n 0.370389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_949_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_950_n 0.0155699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_951_n 0.00601668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_137_74#_c_1029_n 0.00685031f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_62 VNB N_A_593_74#_c_1042_n 0.00204804f $X=-0.19 $Y=-0.245 $X2=1.885
+ $Y2=1.885
cc_63 VNB N_A_593_74#_c_1043_n 0.00204804f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_64 VNB N_A_981_74#_c_1068_n 0.00284399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_981_74#_c_1069_n 0.00215161f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_66 VPB N_C2_c_126_n 0.00832475f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.795
cc_67 VPB N_C2_c_136_n 0.025066f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_68 VPB N_C2_c_137_n 0.0174679f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=1.885
cc_69 VPB N_C2_c_129_n 0.020058f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.635
cc_70 VPB N_C2_c_139_n 0.0205246f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.75
cc_71 VPB N_C2_c_140_n 0.00387294f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.75
cc_72 VPB N_C1_c_225_n 0.0151479f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.495
cc_73 VPB N_C1_c_220_n 0.00324744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_C1_c_221_n 0.00579914f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_75 VPB N_C1_c_228_n 0.0203152f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_76 VPB N_C1_c_229_n 0.0134553f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.75
cc_77 VPB N_B1_c_282_n 0.0387384f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_78 VPB N_B1_c_283_n 0.0348267f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.69
cc_79 VPB N_B1_c_285_n 9.55489e-19 $X=-0.19 $Y=1.66 $X2=1.9 $Y2=0.69
cc_80 VPB N_B1_c_291_n 0.00269836f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_81 VPB N_B1_c_292_n 0.0101177f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.13
cc_82 VPB N_B1_c_293_n 0.00333927f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.665
cc_83 VPB N_B1_c_286_n 0.00184657f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_84 VPB N_B1_c_287_n 0.00153498f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.165
cc_85 VPB N_B2_c_376_n 0.00681642f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.165
cc_86 VPB N_B2_c_382_n 0.0207893f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.69
cc_87 VPB N_B2_c_377_n 0.00705177f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_88 VPB N_B2_c_384_n 0.0222228f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_89 VPB N_B2_c_379_n 0.00323444f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_90 VPB N_A1_c_442_n 0.0332029f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_91 VPB N_A1_c_444_n 0.0423783f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_92 VPB N_A1_c_449_n 0.003453f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_93 VPB N_A1_c_450_n 0.00467714f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.13
cc_94 VPB N_A1_c_451_n 0.00355293f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.665
cc_95 VPB N_A1_c_445_n 0.00180389f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_96 VPB N_A1_c_446_n 0.007317f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.33
cc_97 VPB N_A2_c_532_n 0.0152564f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.495
cc_98 VPB N_A2_c_533_n 0.0150347f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.69
cc_99 VPB A2 0.00212399f $X=-0.19 $Y=1.66 $X2=1.9 $Y2=0.69
cc_100 VPB N_A2_c_531_n 0.0329993f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.75
cc_101 VPB N_Y_c_584_n 0.012628f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.665
cc_102 VPB N_Y_c_586_n 0.0074464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_Y_c_595_n 0.0106598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB Y 0.0155418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB Y 0.0335007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_116_392#_c_732_n 0.00234963f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.13
cc_107 VPB N_A_116_392#_c_733_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.635
cc_108 VPB N_A_116_392#_c_734_n 0.00587129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_116_392#_c_735_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_116_392#_c_736_n 0.0146087f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.33
cc_111 VPB N_A_116_392#_c_737_n 0.00217178f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.33
cc_112 VPB N_A_515_392#_c_791_n 0.00417584f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_113 VPB N_A_515_392#_c_792_n 0.0023327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_515_392#_c_793_n 0.0170232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_515_392#_c_794_n 0.00219816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_515_392#_c_795_n 0.029937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_870_n 0.00329267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_871_n 0.00329129f $X=-0.19 $Y=1.66 $X2=1.9 $Y2=1.13
cc_119 VPB N_VPWR_c_872_n 0.119365f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.13
cc_120 VPB N_VPWR_c_873_n 0.0159778f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_121 VPB N_VPWR_c_874_n 0.0177874f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.33
cc_122 VPB N_VPWR_c_869_n 0.0796337f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.33
cc_123 VPB N_VPWR_c_876_n 0.00656574f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_124 VPB N_VPWR_c_877_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.33
cc_125 N_C2_c_136_n N_C1_c_225_n 0.0205868f $X=0.505 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_126 N_C2_M1014_g N_C1_M1002_g 0.0276308f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_127 N_C2_c_126_n N_C1_c_220_n 0.0058994f $X=0.505 $Y=1.795 $X2=0 $Y2=0
cc_128 N_C2_c_130_n N_C1_c_220_n 0.00312674f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_129 N_C2_c_139_n N_C1_c_220_n 0.00520968f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_130 N_C2_c_129_n N_C1_c_221_n 0.01918f $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_131 N_C2_c_139_n N_C1_c_221_n 0.0117089f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_132 N_C2_c_131_n N_C1_c_221_n 0.00108316f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_133 N_C2_c_137_n N_C1_c_228_n 0.0210693f $X=1.885 $Y=1.885 $X2=0 $Y2=0
cc_134 N_C2_c_139_n N_C1_c_228_n 0.00373749f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_135 N_C2_c_128_n N_C1_M1017_g 0.0224f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_136 N_C2_c_131_n N_C1_M1017_g 0.00174486f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_137 N_C2_c_132_n N_C1_M1017_g 0.00978324f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_138 N_C2_c_126_n N_C1_c_229_n 0.00682553f $X=0.505 $Y=1.795 $X2=0 $Y2=0
cc_139 N_C2_c_139_n N_C1_c_229_n 0.00849886f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_140 N_C2_c_139_n C1 0.0243679f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_141 N_C2_c_131_n C1 0.0110236f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_142 N_C2_c_132_n C1 8.95767e-19 $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_143 C2 C1 0.0265726f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_144 N_C2_c_134_n C1 3.29091e-19 $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_145 N_C2_c_129_n N_C1_c_224_n 0.00978324f $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_146 N_C2_c_139_n N_C1_c_224_n 0.0011826f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_147 C2 N_C1_c_224_n 0.00312674f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_148 N_C2_c_134_n N_C1_c_224_n 0.0213924f $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_149 N_C2_c_132_n N_B1_M1022_g 0.00335539f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_150 N_C2_c_129_n N_B1_c_282_n 0.00519886f $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_151 N_C2_c_136_n N_Y_c_584_n 0.00115778f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_152 N_C2_M1014_g N_Y_c_584_n 0.00514335f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_153 N_C2_c_130_n N_Y_c_584_n 0.00787536f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_154 N_C2_c_140_n N_Y_c_584_n 0.00866338f $X=0.835 $Y=1.75 $X2=0 $Y2=0
cc_155 C2 N_Y_c_584_n 0.0252195f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_156 N_C2_c_134_n N_Y_c_584_n 0.016769f $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_157 N_C2_c_136_n N_Y_c_604_n 0.0143204f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_158 N_C2_c_139_n N_Y_c_604_n 0.0129195f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_159 N_C2_c_140_n N_Y_c_604_n 0.0173978f $X=0.835 $Y=1.75 $X2=0 $Y2=0
cc_160 C2 N_Y_c_604_n 0.00480907f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_161 N_C2_c_134_n N_Y_c_604_n 4.67869e-19 $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_162 N_C2_c_137_n N_Y_c_609_n 0.0164927f $X=1.885 $Y=1.885 $X2=0 $Y2=0
cc_163 N_C2_c_139_n N_Y_c_609_n 0.0424133f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_164 N_C2_c_137_n N_Y_c_586_n 0.00341758f $X=1.885 $Y=1.885 $X2=0 $Y2=0
cc_165 N_C2_c_129_n N_Y_c_586_n 0.00580365f $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_166 N_C2_c_139_n N_Y_c_586_n 0.0137446f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_167 N_C2_c_131_n N_Y_c_586_n 0.0273195f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_168 N_C2_c_128_n N_Y_c_587_n 0.00103145f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_169 N_C2_c_128_n N_Y_c_589_n 0.00440566f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_170 N_C2_c_131_n N_Y_c_589_n 0.0140395f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_171 N_C2_c_132_n N_Y_c_589_n 0.00192034f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_172 N_C2_c_139_n N_Y_c_619_n 0.0193366f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_173 N_C2_M1014_g N_Y_c_620_n 2.14939e-19 $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_174 N_C2_c_128_n N_Y_c_620_n 4.40457e-19 $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_175 N_C2_M1014_g N_Y_c_622_n 0.0133138f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_176 N_C2_c_139_n N_Y_c_622_n 0.00497809f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_177 C2 N_Y_c_622_n 0.0270966f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_178 N_C2_c_134_n N_Y_c_622_n 0.00145942f $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_179 N_C2_c_129_n N_Y_c_595_n 8.62874e-19 $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_180 N_C2_c_139_n N_Y_c_595_n 0.0109918f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_181 N_C2_c_136_n Y 0.00261748f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_182 N_C2_c_136_n Y 0.00631032f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_183 N_C2_c_136_n N_A_116_392#_c_738_n 0.0063803f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_184 N_C2_c_136_n N_A_116_392#_c_733_n 0.00669783f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_C2_c_137_n N_A_116_392#_c_740_n 0.0114481f $X=1.885 $Y=1.885 $X2=0
+ $Y2=0
cc_186 N_C2_c_137_n N_A_116_392#_c_735_n 0.00171731f $X=1.885 $Y=1.885 $X2=0
+ $Y2=0
cc_187 N_C2_c_137_n N_A_116_392#_c_736_n 0.012762f $X=1.885 $Y=1.885 $X2=0 $Y2=0
cc_188 N_C2_c_137_n N_A_515_392#_c_796_n 5.97789e-19 $X=1.885 $Y=1.885 $X2=0
+ $Y2=0
cc_189 N_C2_c_136_n N_VPWR_c_872_n 0.0044313f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_190 N_C2_c_137_n N_VPWR_c_872_n 0.00278257f $X=1.885 $Y=1.885 $X2=0 $Y2=0
cc_191 N_C2_c_136_n N_VPWR_c_869_n 0.00857701f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_192 N_C2_c_137_n N_VPWR_c_869_n 0.00358707f $X=1.885 $Y=1.885 $X2=0 $Y2=0
cc_193 N_C2_M1014_g N_VGND_c_941_n 0.0105743f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_194 N_C2_c_128_n N_VGND_c_942_n 0.0118294f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_195 N_C2_c_131_n N_VGND_c_942_n 0.0114324f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_196 N_C2_c_132_n N_VGND_c_942_n 9.66467e-19 $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_197 N_C2_M1014_g N_VGND_c_944_n 0.00433162f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_198 N_C2_c_128_n N_VGND_c_944_n 0.00383152f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_199 N_C2_M1014_g N_VGND_c_948_n 0.00446997f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_200 N_C2_c_128_n N_VGND_c_948_n 0.00757637f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_201 N_C2_M1014_g N_A_137_74#_c_1029_n 0.00366414f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_202 N_C2_c_128_n N_A_137_74#_c_1029_n 7.20798e-19 $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_203 N_C1_c_225_n N_Y_c_604_n 0.0126342f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_204 N_C1_c_228_n N_Y_c_609_n 0.0126342f $X=1.435 $Y=1.885 $X2=0 $Y2=0
cc_205 N_C1_c_229_n N_Y_c_619_n 0.00137147f $X=1.04 $Y=1.81 $X2=0 $Y2=0
cc_206 N_C1_M1002_g N_Y_c_620_n 0.00185091f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_207 N_C1_M1017_g N_Y_c_620_n 0.00411699f $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_208 N_C1_c_224_n N_Y_c_620_n 7.12379e-19 $X=1.47 $Y=1.33 $X2=0 $Y2=0
cc_209 N_C1_M1002_g N_Y_c_622_n 0.00815093f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_210 C1 N_Y_c_622_n 0.0221715f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_211 N_C1_c_225_n N_A_116_392#_c_738_n 0.00714743f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_212 N_C1_c_228_n N_A_116_392#_c_738_n 5.36851e-19 $X=1.435 $Y=1.885 $X2=0
+ $Y2=0
cc_213 N_C1_c_225_n N_A_116_392#_c_732_n 0.0110098f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_214 N_C1_c_228_n N_A_116_392#_c_732_n 0.0110098f $X=1.435 $Y=1.885 $X2=0
+ $Y2=0
cc_215 N_C1_c_225_n N_A_116_392#_c_733_n 0.00171731f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_C1_c_225_n N_A_116_392#_c_740_n 5.36851e-19 $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_C1_c_228_n N_A_116_392#_c_740_n 0.00714743f $X=1.435 $Y=1.885 $X2=0
+ $Y2=0
cc_218 N_C1_c_228_n N_A_116_392#_c_735_n 0.00171731f $X=1.435 $Y=1.885 $X2=0
+ $Y2=0
cc_219 N_C1_c_225_n N_VPWR_c_872_n 0.00278257f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_220 N_C1_c_228_n N_VPWR_c_872_n 0.00278257f $X=1.435 $Y=1.885 $X2=0 $Y2=0
cc_221 N_C1_c_225_n N_VPWR_c_869_n 0.00354187f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_222 N_C1_c_228_n N_VPWR_c_869_n 0.00354187f $X=1.435 $Y=1.885 $X2=0 $Y2=0
cc_223 N_C1_M1017_g N_VGND_c_942_n 9.22378e-19 $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_224 N_C1_M1002_g N_VGND_c_944_n 0.00291649f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_225 N_C1_M1017_g N_VGND_c_944_n 0.00291649f $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_226 N_C1_M1002_g N_VGND_c_948_n 0.00359219f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_227 N_C1_M1017_g N_VGND_c_948_n 0.00359219f $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_228 N_C1_M1002_g N_A_137_74#_c_1029_n 0.0106323f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_229 N_C1_M1017_g N_A_137_74#_c_1029_n 0.0156912f $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_230 N_B1_M1022_g N_B2_M1015_g 0.040022f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_231 N_B1_c_282_n N_B2_c_376_n 0.0121603f $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_232 N_B1_c_285_n N_B2_c_376_n 0.00204043f $X=3.15 $Y=1.8 $X2=0 $Y2=0
cc_233 N_B1_c_282_n N_B2_c_382_n 0.0345528f $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_234 N_B1_c_291_n N_B2_c_382_n 0.00346066f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_235 N_B1_c_292_n N_B2_c_382_n 0.0140592f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_236 N_B1_c_283_n N_B2_c_377_n 0.00263656f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_237 N_B1_c_293_n N_B2_c_377_n 0.00227237f $X=4.19 $Y=1.95 $X2=0 $Y2=0
cc_238 N_B1_c_283_n N_B2_c_384_n 0.0260686f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_239 N_B1_c_292_n N_B2_c_384_n 0.0167929f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_240 N_B1_c_293_n N_B2_c_384_n 0.0013695f $X=4.19 $Y=1.95 $X2=0 $Y2=0
cc_241 N_B1_M1023_g N_B2_c_378_n 0.0286129f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_242 N_B1_M1022_g N_B2_c_379_n 8.86752e-19 $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_243 N_B1_c_282_n N_B2_c_379_n 2.29946e-19 $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_244 N_B1_M1023_g N_B2_c_379_n 7.75734e-19 $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_245 N_B1_c_285_n N_B2_c_379_n 0.0256873f $X=3.15 $Y=1.8 $X2=0 $Y2=0
cc_246 N_B1_c_292_n N_B2_c_379_n 0.0265118f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_247 N_B1_c_286_n N_B2_c_379_n 0.0154943f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_248 N_B1_c_282_n N_B2_c_380_n 0.00781816f $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_249 N_B1_c_283_n N_B2_c_380_n 0.0206191f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_250 N_B1_M1023_g N_B2_c_380_n 0.00771183f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_251 N_B1_c_285_n N_B2_c_380_n 0.00109171f $X=3.15 $Y=1.8 $X2=0 $Y2=0
cc_252 N_B1_c_292_n N_B2_c_380_n 0.00243942f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_253 N_B1_c_286_n N_B2_c_380_n 0.00273929f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_254 N_B1_M1023_g N_A1_M1011_g 0.0266162f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_255 N_B1_c_283_n N_A1_c_442_n 0.0343429f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_256 N_B1_c_286_n N_A1_c_442_n 4.14342e-19 $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_257 N_B1_c_293_n N_A1_c_449_n 0.00477463f $X=4.19 $Y=1.95 $X2=0 $Y2=0
cc_258 N_B1_c_283_n N_A1_c_445_n 4.13565e-19 $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_259 N_B1_c_286_n N_A1_c_445_n 0.0215802f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_260 N_B1_M1022_g N_Y_c_586_n 0.00329148f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_261 N_B1_c_282_n N_Y_c_586_n 0.00423475f $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_262 N_B1_c_291_n N_Y_c_586_n 0.00462099f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_263 N_B1_c_331_p N_Y_c_586_n 4.83905e-19 $X=3.235 $Y=2.035 $X2=0 $Y2=0
cc_264 N_B1_c_287_n N_Y_c_586_n 0.0219971f $X=3.065 $Y=1.635 $X2=0 $Y2=0
cc_265 N_B1_M1022_g N_Y_c_587_n 0.0078351f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_266 N_B1_M1022_g N_Y_c_588_n 0.0120432f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_267 N_B1_c_282_n N_Y_c_588_n 0.00153394f $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_268 N_B1_c_283_n N_Y_c_588_n 0.00358406f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_269 N_B1_M1023_g N_Y_c_588_n 0.0197687f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_270 N_B1_c_285_n N_Y_c_588_n 0.00818622f $X=3.15 $Y=1.8 $X2=0 $Y2=0
cc_271 N_B1_c_286_n N_Y_c_588_n 0.0164207f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_272 N_B1_c_287_n N_Y_c_588_n 0.00888366f $X=3.065 $Y=1.635 $X2=0 $Y2=0
cc_273 N_B1_M1022_g N_Y_c_589_n 0.0104367f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_274 N_B1_c_282_n N_Y_c_589_n 0.00326139f $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_275 N_B1_c_287_n N_Y_c_589_n 0.0138023f $X=3.065 $Y=1.635 $X2=0 $Y2=0
cc_276 N_B1_M1023_g N_Y_c_590_n 0.00756015f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_277 N_B1_c_282_n N_Y_c_595_n 4.21939e-19 $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_278 N_B1_c_292_n N_A_116_392#_M1005_s 2.87715e-19 $X=4.105 $Y=2.035 $X2=0
+ $Y2=0
cc_279 N_B1_c_331_p N_A_116_392#_M1005_s 0.00221065f $X=3.235 $Y=2.035 $X2=0
+ $Y2=0
cc_280 N_B1_c_292_n N_A_116_392#_M1021_s 0.00423457f $X=4.105 $Y=2.035 $X2=0
+ $Y2=0
cc_281 N_B1_c_283_n N_A_116_392#_c_734_n 0.00378312f $X=4.385 $Y=1.885 $X2=0
+ $Y2=0
cc_282 N_B1_c_282_n N_A_116_392#_c_736_n 0.00994772f $X=2.945 $Y=1.885 $X2=0
+ $Y2=0
cc_283 N_B1_c_282_n N_A_116_392#_c_737_n 0.0108919f $X=2.945 $Y=1.885 $X2=0
+ $Y2=0
cc_284 N_B1_c_292_n N_A_515_392#_M1020_d 0.00198204f $X=4.105 $Y=2.035 $X2=0
+ $Y2=0
cc_285 N_B1_c_282_n N_A_515_392#_c_796_n 0.00300514f $X=2.945 $Y=1.885 $X2=0
+ $Y2=0
cc_286 N_B1_c_287_n N_A_515_392#_c_796_n 0.0106529f $X=3.065 $Y=1.635 $X2=0
+ $Y2=0
cc_287 N_B1_c_282_n N_A_515_392#_c_800_n 0.0131184f $X=2.945 $Y=1.885 $X2=0
+ $Y2=0
cc_288 N_B1_c_283_n N_A_515_392#_c_800_n 0.0137087f $X=4.385 $Y=1.885 $X2=0
+ $Y2=0
cc_289 N_B1_c_292_n N_A_515_392#_c_800_n 0.0564308f $X=4.105 $Y=2.035 $X2=0
+ $Y2=0
cc_290 N_B1_c_331_p N_A_515_392#_c_800_n 0.0128074f $X=3.235 $Y=2.035 $X2=0
+ $Y2=0
cc_291 N_B1_c_286_n N_A_515_392#_c_800_n 0.004488f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_292 N_B1_c_287_n N_A_515_392#_c_800_n 0.00647386f $X=3.065 $Y=1.635 $X2=0
+ $Y2=0
cc_293 N_B1_c_283_n N_A_515_392#_c_791_n 0.0056206f $X=4.385 $Y=1.885 $X2=0
+ $Y2=0
cc_294 N_B1_c_292_n N_A_515_392#_c_791_n 0.00682867f $X=4.105 $Y=2.035 $X2=0
+ $Y2=0
cc_295 N_B1_c_286_n N_A_515_392#_c_791_n 0.00232751f $X=4.31 $Y=1.615 $X2=0
+ $Y2=0
cc_296 N_B1_c_283_n N_A_515_392#_c_794_n 8.50317e-19 $X=4.385 $Y=1.885 $X2=0
+ $Y2=0
cc_297 N_B1_c_283_n N_VPWR_c_870_n 6.25687e-19 $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_298 N_B1_c_282_n N_VPWR_c_872_n 0.00278271f $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_299 N_B1_c_283_n N_VPWR_c_872_n 0.00444483f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_300 N_B1_c_282_n N_VPWR_c_869_n 0.00358708f $X=2.945 $Y=1.885 $X2=0 $Y2=0
cc_301 N_B1_c_283_n N_VPWR_c_869_n 0.00855608f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_302 N_B1_M1022_g N_VGND_c_942_n 0.00380203f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_303 N_B1_M1022_g N_VGND_c_945_n 0.00434272f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_304 N_B1_M1023_g N_VGND_c_946_n 0.00434272f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_305 N_B1_M1022_g N_VGND_c_948_n 0.00826366f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_306 N_B1_M1023_g N_VGND_c_948_n 0.00821465f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_307 N_B2_M1015_g N_Y_c_587_n 9.56968e-19 $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_308 N_B2_M1015_g N_Y_c_588_n 0.0158888f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_309 N_B2_c_378_n N_Y_c_588_n 0.0153959f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_310 N_B2_c_379_n N_Y_c_588_n 0.0256597f $X=3.57 $Y=1.425 $X2=0 $Y2=0
cc_311 N_B2_c_380_n N_Y_c_588_n 0.0113378f $X=3.845 $Y=1.34 $X2=0 $Y2=0
cc_312 N_B2_M1015_g N_Y_c_589_n 9.79153e-19 $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_313 N_B2_c_379_n N_Y_c_589_n 0.00116356f $X=3.57 $Y=1.425 $X2=0 $Y2=0
cc_314 N_B2_c_378_n N_Y_c_590_n 9.65066e-19 $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_315 N_B2_c_382_n N_A_116_392#_c_734_n 0.0116178f $X=3.395 $Y=1.885 $X2=0
+ $Y2=0
cc_316 N_B2_c_384_n N_A_116_392#_c_734_n 0.0127359f $X=3.845 $Y=1.885 $X2=0
+ $Y2=0
cc_317 N_B2_c_382_n N_A_116_392#_c_737_n 0.00427652f $X=3.395 $Y=1.885 $X2=0
+ $Y2=0
cc_318 N_B2_c_384_n N_A_116_392#_c_737_n 5.32705e-19 $X=3.845 $Y=1.885 $X2=0
+ $Y2=0
cc_319 N_B2_c_382_n N_A_515_392#_c_800_n 0.00862059f $X=3.395 $Y=1.885 $X2=0
+ $Y2=0
cc_320 N_B2_c_384_n N_A_515_392#_c_800_n 0.00908392f $X=3.845 $Y=1.885 $X2=0
+ $Y2=0
cc_321 N_B2_c_384_n N_A_515_392#_c_791_n 8.86046e-19 $X=3.845 $Y=1.885 $X2=0
+ $Y2=0
cc_322 N_B2_c_382_n N_VPWR_c_872_n 0.00290311f $X=3.395 $Y=1.885 $X2=0 $Y2=0
cc_323 N_B2_c_384_n N_VPWR_c_872_n 0.00291649f $X=3.845 $Y=1.885 $X2=0 $Y2=0
cc_324 N_B2_c_382_n N_VPWR_c_869_n 0.0035903f $X=3.395 $Y=1.885 $X2=0 $Y2=0
cc_325 N_B2_c_384_n N_VPWR_c_869_n 0.00360347f $X=3.845 $Y=1.885 $X2=0 $Y2=0
cc_326 N_B2_M1015_g N_VGND_c_945_n 0.00316493f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_327 N_B2_c_378_n N_VGND_c_946_n 0.00316493f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_328 N_B2_M1015_g N_VGND_c_948_n 0.00393725f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_329 N_B2_c_378_n N_VGND_c_948_n 0.00393725f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_330 N_B2_M1015_g N_VGND_c_950_n 0.00381881f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_331 N_B2_c_378_n N_VGND_c_950_n 0.00381881f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_332 N_B2_M1015_g N_A_593_74#_c_1044_n 0.00966972f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_333 N_B2_c_378_n N_A_593_74#_c_1044_n 0.00966972f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_334 N_B2_M1015_g N_A_593_74#_c_1042_n 0.00590335f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_335 N_B2_c_378_n N_A_593_74#_c_1042_n 8.35363e-19 $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_336 N_B2_M1015_g N_A_593_74#_c_1043_n 8.35363e-19 $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_337 N_B2_c_378_n N_A_593_74#_c_1043_n 0.00590335f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_338 N_A1_c_442_n N_A2_c_532_n 0.0285051f $X=4.835 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_339 N_A1_c_449_n N_A2_c_532_n 0.0014352f $X=5.03 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_340 N_A1_c_450_n N_A2_c_532_n 0.0114321f $X=5.885 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_341 N_A1_M1011_g N_A2_M1000_g 0.0300052f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_342 N_A1_c_444_n N_A2_c_533_n 0.0321416f $X=6.215 $Y=1.885 $X2=0 $Y2=0
cc_343 N_A1_c_450_n N_A2_c_533_n 0.0124528f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_344 N_A1_c_451_n N_A2_c_533_n 0.00156409f $X=5.97 $Y=1.95 $X2=0 $Y2=0
cc_345 N_A1_M1013_g N_A2_M1001_g 0.0266095f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_346 N_A1_c_442_n A2 2.99931e-19 $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_347 N_A1_c_444_n A2 2.19852e-19 $X=6.215 $Y=1.885 $X2=0 $Y2=0
cc_348 N_A1_c_450_n A2 0.0244586f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_349 N_A1_c_445_n A2 0.0244979f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_350 N_A1_c_446_n A2 0.0204271f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_351 N_A1_c_442_n N_A2_c_531_n 0.0249247f $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_352 N_A1_c_444_n N_A2_c_531_n 0.0193662f $X=6.215 $Y=1.885 $X2=0 $Y2=0
cc_353 N_A1_c_449_n N_A2_c_531_n 0.00238087f $X=5.03 $Y=1.95 $X2=0 $Y2=0
cc_354 N_A1_c_450_n N_A2_c_531_n 0.00486801f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_355 N_A1_c_451_n N_A2_c_531_n 0.00259167f $X=5.97 $Y=1.95 $X2=0 $Y2=0
cc_356 N_A1_c_445_n N_A2_c_531_n 0.00243494f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_357 N_A1_c_446_n N_A2_c_531_n 0.00375221f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_358 N_A1_M1011_g N_Y_c_588_n 3.91998e-19 $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_359 N_A1_c_442_n N_Y_c_588_n 6.75574e-19 $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_360 N_A1_c_445_n N_Y_c_588_n 0.00244567f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_361 N_A1_M1011_g N_Y_c_590_n 0.00279931f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_362 N_A1_M1011_g N_Y_c_591_n 0.0135003f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_363 N_A1_c_442_n N_Y_c_591_n 0.00341567f $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_364 N_A1_M1013_g N_Y_c_591_n 0.0156502f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_365 N_A1_c_444_n N_Y_c_591_n 0.00423048f $X=6.215 $Y=1.885 $X2=0 $Y2=0
cc_366 N_A1_c_450_n N_Y_c_591_n 0.0111742f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_367 N_A1_c_445_n N_Y_c_591_n 0.0299139f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_368 N_A1_c_446_n N_Y_c_591_n 0.0444698f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_369 N_A1_M1013_g N_Y_c_592_n 0.00453147f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_370 N_A1_c_450_n N_A_515_392#_M1003_d 0.00197722f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_371 N_A1_c_442_n N_A_515_392#_c_791_n 0.00681585f $X=4.835 $Y=1.885 $X2=0
+ $Y2=0
cc_372 N_A1_c_494_p N_A_515_392#_c_791_n 0.00682867f $X=5.115 $Y=2.035 $X2=0
+ $Y2=0
cc_373 N_A1_c_445_n N_A_515_392#_c_791_n 0.00734325f $X=5.03 $Y=1.615 $X2=0
+ $Y2=0
cc_374 N_A1_c_442_n N_A_515_392#_c_817_n 0.0114849f $X=4.835 $Y=1.885 $X2=0
+ $Y2=0
cc_375 N_A1_c_450_n N_A_515_392#_c_817_n 0.0151646f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_376 N_A1_c_494_p N_A_515_392#_c_817_n 0.0114873f $X=5.115 $Y=2.035 $X2=0
+ $Y2=0
cc_377 N_A1_c_445_n N_A_515_392#_c_817_n 0.00451997f $X=5.03 $Y=1.615 $X2=0
+ $Y2=0
cc_378 N_A1_c_444_n N_A_515_392#_c_821_n 0.0110913f $X=6.215 $Y=1.885 $X2=0
+ $Y2=0
cc_379 N_A1_c_450_n N_A_515_392#_c_821_n 0.0224835f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_380 N_A1_c_446_n N_A_515_392#_c_821_n 0.00603861f $X=6.29 $Y=1.615 $X2=0
+ $Y2=0
cc_381 N_A1_c_444_n N_A_515_392#_c_793_n 0.00908089f $X=6.215 $Y=1.885 $X2=0
+ $Y2=0
cc_382 N_A1_c_450_n N_A_515_392#_c_793_n 0.0115259f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_383 N_A1_c_446_n N_A_515_392#_c_793_n 0.0149332f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_384 N_A1_c_442_n N_A_515_392#_c_794_n 5.94216e-19 $X=4.835 $Y=1.885 $X2=0
+ $Y2=0
cc_385 N_A1_c_450_n N_A_515_392#_c_828_n 0.0151508f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_386 N_A1_c_444_n N_A_515_392#_c_795_n 0.00149863f $X=6.215 $Y=1.885 $X2=0
+ $Y2=0
cc_387 N_A1_c_450_n N_VPWR_M1006_s 7.13959e-19 $X=5.885 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_388 N_A1_c_494_p N_VPWR_M1006_s 0.0023739f $X=5.115 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_389 N_A1_c_450_n N_VPWR_M1004_s 0.00350478f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_390 N_A1_c_442_n N_VPWR_c_870_n 0.00737663f $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_391 N_A1_c_444_n N_VPWR_c_871_n 0.00937738f $X=6.215 $Y=1.885 $X2=0 $Y2=0
cc_392 N_A1_c_442_n N_VPWR_c_872_n 0.00413917f $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_393 N_A1_c_444_n N_VPWR_c_874_n 0.00413917f $X=6.215 $Y=1.885 $X2=0 $Y2=0
cc_394 N_A1_c_442_n N_VPWR_c_869_n 0.00416821f $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_395 N_A1_c_444_n N_VPWR_c_869_n 0.00420231f $X=6.215 $Y=1.885 $X2=0 $Y2=0
cc_396 N_A1_M1011_g N_VGND_c_943_n 5.94048e-19 $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_397 N_A1_M1013_g N_VGND_c_943_n 5.48301e-19 $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_398 N_A1_M1011_g N_VGND_c_946_n 0.00439937f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_399 N_A1_M1013_g N_VGND_c_947_n 0.00433834f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_400 N_A1_M1011_g N_VGND_c_948_n 0.00840422f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_401 N_A1_M1013_g N_VGND_c_948_n 0.00824802f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_402 N_A1_M1011_g N_A_981_74#_c_1068_n 0.00450875f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_403 N_A1_M1011_g N_A_981_74#_c_1071_n 0.00192658f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_404 N_A1_M1013_g N_A_981_74#_c_1072_n 0.00215008f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_405 N_A1_M1013_g N_A_981_74#_c_1069_n 0.00587363f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_406 N_A2_M1000_g N_Y_c_591_n 0.011602f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_407 N_A2_M1001_g N_Y_c_591_n 0.0127746f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_408 A2 N_Y_c_591_n 0.0244045f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_409 N_A2_c_531_n N_Y_c_591_n 0.00196123f $X=5.765 $Y=1.667 $X2=0 $Y2=0
cc_410 N_A2_c_532_n N_A_515_392#_c_791_n 9.12982e-19 $X=5.315 $Y=1.885 $X2=0
+ $Y2=0
cc_411 N_A2_c_532_n N_A_515_392#_c_817_n 0.0105707f $X=5.315 $Y=1.885 $X2=0
+ $Y2=0
cc_412 N_A2_c_532_n N_A_515_392#_c_792_n 3.38692e-19 $X=5.315 $Y=1.885 $X2=0
+ $Y2=0
cc_413 N_A2_c_533_n N_A_515_392#_c_792_n 3.38692e-19 $X=5.765 $Y=1.885 $X2=0
+ $Y2=0
cc_414 N_A2_c_533_n N_A_515_392#_c_821_n 0.0103891f $X=5.765 $Y=1.885 $X2=0
+ $Y2=0
cc_415 N_A2_c_533_n N_A_515_392#_c_793_n 9.37611e-19 $X=5.765 $Y=1.885 $X2=0
+ $Y2=0
cc_416 N_A2_c_532_n N_VPWR_c_870_n 0.00722898f $X=5.315 $Y=1.885 $X2=0 $Y2=0
cc_417 N_A2_c_533_n N_VPWR_c_870_n 4.12151e-19 $X=5.765 $Y=1.885 $X2=0 $Y2=0
cc_418 N_A2_c_532_n N_VPWR_c_871_n 4.12446e-19 $X=5.315 $Y=1.885 $X2=0 $Y2=0
cc_419 N_A2_c_533_n N_VPWR_c_871_n 0.00710435f $X=5.765 $Y=1.885 $X2=0 $Y2=0
cc_420 N_A2_c_532_n N_VPWR_c_873_n 0.00413917f $X=5.315 $Y=1.885 $X2=0 $Y2=0
cc_421 N_A2_c_533_n N_VPWR_c_873_n 0.00413917f $X=5.765 $Y=1.885 $X2=0 $Y2=0
cc_422 N_A2_c_532_n N_VPWR_c_869_n 0.00416762f $X=5.315 $Y=1.885 $X2=0 $Y2=0
cc_423 N_A2_c_533_n N_VPWR_c_869_n 0.00416762f $X=5.765 $Y=1.885 $X2=0 $Y2=0
cc_424 N_A2_M1000_g N_VGND_c_943_n 0.00681232f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_425 N_A2_M1001_g N_VGND_c_943_n 0.0066056f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_426 N_A2_M1000_g N_VGND_c_946_n 0.00398535f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_427 N_A2_M1001_g N_VGND_c_947_n 0.00398535f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_428 N_A2_M1000_g N_VGND_c_948_n 0.00384569f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_429 N_A2_M1001_g N_VGND_c_948_n 0.00383955f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_430 N_A2_M1000_g N_A_981_74#_c_1068_n 0.00227555f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_431 N_A2_M1000_g N_A_981_74#_c_1075_n 0.0119053f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_432 N_A2_M1001_g N_A_981_74#_c_1075_n 0.00951514f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_433 N_A2_M1001_g N_A_981_74#_c_1069_n 2.96277e-19 $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_434 N_Y_c_604_n N_A_116_392#_M1009_d 0.00381853f $X=1.065 $Y=2.09 $X2=-0.19
+ $Y2=-0.245
cc_435 N_Y_c_609_n N_A_116_392#_M1010_d 0.00395925f $X=1.995 $Y=2.09 $X2=0 $Y2=0
cc_436 N_Y_c_604_n N_A_116_392#_c_738_n 0.0171814f $X=1.065 $Y=2.09 $X2=0 $Y2=0
cc_437 Y N_A_116_392#_c_738_n 0.0378419f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_438 N_Y_M1007_s N_A_116_392#_c_732_n 0.00229612f $X=1.03 $Y=1.96 $X2=0 $Y2=0
cc_439 N_Y_c_685_p N_A_116_392#_c_732_n 0.0164404f $X=1.195 $Y=2.57 $X2=0 $Y2=0
cc_440 Y N_A_116_392#_c_733_n 0.00541333f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_441 N_Y_c_609_n N_A_116_392#_c_740_n 0.0171814f $X=1.995 $Y=2.09 $X2=0 $Y2=0
cc_442 N_Y_M1012_s N_A_116_392#_c_736_n 0.00355467f $X=1.96 $Y=1.96 $X2=0 $Y2=0
cc_443 N_Y_c_595_n N_A_116_392#_c_736_n 0.0344828f $X=2.16 $Y=2.17 $X2=0 $Y2=0
cc_444 N_Y_c_586_n N_A_515_392#_c_796_n 0.00255114f $X=2.38 $Y=2.005 $X2=0 $Y2=0
cc_445 N_Y_c_589_n N_A_515_392#_c_796_n 0.0013185f $X=2.84 $Y=1.005 $X2=0 $Y2=0
cc_446 N_Y_c_595_n N_A_515_392#_c_796_n 0.0232784f $X=2.16 $Y=2.17 $X2=0 $Y2=0
cc_447 N_Y_c_595_n N_A_515_392#_c_839_n 0.0220283f $X=2.16 $Y=2.17 $X2=0 $Y2=0
cc_448 N_Y_c_588_n N_A_515_392#_c_791_n 0.00748381f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_449 N_Y_c_591_n N_A_515_392#_c_793_n 0.0044659f $X=6.32 $Y=1.195 $X2=0 $Y2=0
cc_450 N_Y_c_595_n N_A_515_392#_c_842_n 0.0151273f $X=2.16 $Y=2.17 $X2=0 $Y2=0
cc_451 Y N_VPWR_c_872_n 0.0124046f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_452 Y N_VPWR_c_869_n 0.0102675f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_453 N_Y_c_584_n N_VGND_M1014_d 2.6293e-19 $X=0.17 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_454 N_Y_c_585_n N_VGND_M1014_d 0.00243255f $X=0.255 $Y=0.91 $X2=-0.19
+ $Y2=-0.245
cc_455 N_Y_c_622_n N_VGND_M1014_d 0.00982502f $X=1.09 $Y=0.887 $X2=-0.19
+ $Y2=-0.245
cc_456 N_Y_c_588_n N_VGND_M1015_d 0.00480292f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_457 N_Y_c_585_n N_VGND_c_941_n 0.0122781f $X=0.255 $Y=0.91 $X2=0 $Y2=0
cc_458 N_Y_c_622_n N_VGND_c_941_n 0.0176875f $X=1.09 $Y=0.887 $X2=0 $Y2=0
cc_459 N_Y_c_587_n N_VGND_c_942_n 0.0383948f $X=2.675 $Y=0.515 $X2=0 $Y2=0
cc_460 N_Y_c_589_n N_VGND_c_942_n 0.00143078f $X=2.84 $Y=1.005 $X2=0 $Y2=0
cc_461 N_Y_c_620_n N_VGND_c_942_n 0.00172463f $X=1.255 $Y=0.865 $X2=0 $Y2=0
cc_462 N_Y_c_587_n N_VGND_c_945_n 0.0145639f $X=2.675 $Y=0.515 $X2=0 $Y2=0
cc_463 N_Y_c_590_n N_VGND_c_946_n 0.0116636f $X=4.615 $Y=0.515 $X2=0 $Y2=0
cc_464 N_Y_c_592_n N_VGND_c_947_n 0.0115122f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_465 N_Y_c_585_n N_VGND_c_948_n 0.00175584f $X=0.255 $Y=0.91 $X2=0 $Y2=0
cc_466 N_Y_c_587_n N_VGND_c_948_n 0.0119984f $X=2.675 $Y=0.515 $X2=0 $Y2=0
cc_467 N_Y_c_590_n N_VGND_c_948_n 0.00959771f $X=4.615 $Y=0.515 $X2=0 $Y2=0
cc_468 N_Y_c_592_n N_VGND_c_948_n 0.0095288f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_469 N_Y_c_622_n N_VGND_c_948_n 0.00688546f $X=1.09 $Y=0.887 $X2=0 $Y2=0
cc_470 N_Y_c_622_n N_A_137_74#_M1014_s 0.00441403f $X=1.09 $Y=0.887 $X2=-0.19
+ $Y2=-0.245
cc_471 N_Y_M1002_s N_A_137_74#_c_1029_n 0.0016448f $X=1.115 $Y=0.37 $X2=0 $Y2=0
cc_472 N_Y_c_620_n N_A_137_74#_c_1029_n 0.0156706f $X=1.255 $Y=0.865 $X2=0 $Y2=0
cc_473 N_Y_c_622_n N_A_137_74#_c_1029_n 0.0181933f $X=1.09 $Y=0.887 $X2=0 $Y2=0
cc_474 N_Y_c_588_n N_A_593_74#_M1022_d 0.00176461f $X=4.45 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_475 N_Y_c_588_n N_A_593_74#_M1018_s 0.00176461f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_476 N_Y_c_588_n N_A_593_74#_c_1044_n 0.0449815f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_477 N_Y_c_587_n N_A_593_74#_c_1042_n 0.0150645f $X=2.675 $Y=0.515 $X2=0 $Y2=0
cc_478 N_Y_c_588_n N_A_593_74#_c_1042_n 0.0146914f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_479 N_Y_c_588_n N_A_593_74#_c_1043_n 0.0146914f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_480 N_Y_c_590_n N_A_593_74#_c_1043_n 0.0145907f $X=4.615 $Y=0.515 $X2=0 $Y2=0
cc_481 N_Y_c_590_n N_A_981_74#_c_1068_n 0.0164865f $X=4.615 $Y=0.515 $X2=0 $Y2=0
cc_482 N_Y_c_591_n N_A_981_74#_c_1075_n 0.0411874f $X=6.32 $Y=1.195 $X2=0 $Y2=0
cc_483 N_Y_c_591_n N_A_981_74#_c_1071_n 0.023557f $X=6.32 $Y=1.195 $X2=0 $Y2=0
cc_484 N_Y_c_591_n N_A_981_74#_c_1072_n 0.0176844f $X=6.32 $Y=1.195 $X2=0 $Y2=0
cc_485 N_Y_c_592_n N_A_981_74#_c_1069_n 0.0158295f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_486 N_A_116_392#_c_736_n N_A_515_392#_M1005_d 0.00459288f $X=3.005 $Y=2.852
+ $X2=-0.19 $Y2=1.66
cc_487 N_A_116_392#_c_734_n N_A_515_392#_M1020_d 0.0021207f $X=4.115 $Y=2.815
+ $X2=0 $Y2=0
cc_488 N_A_116_392#_c_736_n N_A_515_392#_c_839_n 0.012787f $X=3.005 $Y=2.852
+ $X2=0 $Y2=0
cc_489 N_A_116_392#_c_737_n N_A_515_392#_c_839_n 0.00713087f $X=3.335 $Y=2.852
+ $X2=0 $Y2=0
cc_490 N_A_116_392#_M1005_s N_A_515_392#_c_800_n 0.00395998f $X=3.02 $Y=1.96
+ $X2=0 $Y2=0
cc_491 N_A_116_392#_M1021_s N_A_515_392#_c_800_n 0.00617463f $X=3.92 $Y=1.96
+ $X2=0 $Y2=0
cc_492 N_A_116_392#_c_734_n N_A_515_392#_c_800_n 0.0519419f $X=4.115 $Y=2.815
+ $X2=0 $Y2=0
cc_493 N_A_116_392#_c_736_n N_A_515_392#_c_800_n 0.00443481f $X=3.005 $Y=2.852
+ $X2=0 $Y2=0
cc_494 N_A_116_392#_c_737_n N_A_515_392#_c_800_n 0.016671f $X=3.335 $Y=2.852
+ $X2=0 $Y2=0
cc_495 N_A_116_392#_c_734_n N_A_515_392#_c_794_n 0.0141875f $X=4.115 $Y=2.815
+ $X2=0 $Y2=0
cc_496 N_A_116_392#_c_732_n N_VPWR_c_872_n 0.0378125f $X=1.495 $Y=2.99 $X2=0
+ $Y2=0
cc_497 N_A_116_392#_c_733_n N_VPWR_c_872_n 0.0235512f $X=0.895 $Y=2.99 $X2=0
+ $Y2=0
cc_498 N_A_116_392#_c_734_n N_VPWR_c_872_n 0.0409513f $X=4.115 $Y=2.815 $X2=0
+ $Y2=0
cc_499 N_A_116_392#_c_735_n N_VPWR_c_872_n 0.0235512f $X=1.66 $Y=2.99 $X2=0
+ $Y2=0
cc_500 N_A_116_392#_c_736_n N_VPWR_c_872_n 0.0978434f $X=3.005 $Y=2.852 $X2=0
+ $Y2=0
cc_501 N_A_116_392#_c_732_n N_VPWR_c_869_n 0.0213231f $X=1.495 $Y=2.99 $X2=0
+ $Y2=0
cc_502 N_A_116_392#_c_733_n N_VPWR_c_869_n 0.0126924f $X=0.895 $Y=2.99 $X2=0
+ $Y2=0
cc_503 N_A_116_392#_c_734_n N_VPWR_c_869_n 0.0342454f $X=4.115 $Y=2.815 $X2=0
+ $Y2=0
cc_504 N_A_116_392#_c_735_n N_VPWR_c_869_n 0.0126924f $X=1.66 $Y=2.99 $X2=0
+ $Y2=0
cc_505 N_A_116_392#_c_736_n N_VPWR_c_869_n 0.0556764f $X=3.005 $Y=2.852 $X2=0
+ $Y2=0
cc_506 N_A_515_392#_c_817_n N_VPWR_M1006_s 0.00452475f $X=5.425 $Y=2.385
+ $X2=-0.19 $Y2=1.66
cc_507 N_A_515_392#_c_821_n N_VPWR_M1004_s 0.00415698f $X=6.275 $Y=2.385 $X2=0
+ $Y2=0
cc_508 N_A_515_392#_c_817_n N_VPWR_c_870_n 0.0193487f $X=5.425 $Y=2.385 $X2=0
+ $Y2=0
cc_509 N_A_515_392#_c_792_n N_VPWR_c_870_n 0.0132968f $X=5.54 $Y=2.815 $X2=0
+ $Y2=0
cc_510 N_A_515_392#_c_794_n N_VPWR_c_870_n 0.0126977f $X=4.61 $Y=2.465 $X2=0
+ $Y2=0
cc_511 N_A_515_392#_c_792_n N_VPWR_c_871_n 0.0131308f $X=5.54 $Y=2.815 $X2=0
+ $Y2=0
cc_512 N_A_515_392#_c_821_n N_VPWR_c_871_n 0.0169419f $X=6.275 $Y=2.385 $X2=0
+ $Y2=0
cc_513 N_A_515_392#_c_795_n N_VPWR_c_871_n 0.0140562f $X=6.44 $Y=2.455 $X2=0
+ $Y2=0
cc_514 N_A_515_392#_c_794_n N_VPWR_c_872_n 0.00950426f $X=4.61 $Y=2.465 $X2=0
+ $Y2=0
cc_515 N_A_515_392#_c_792_n N_VPWR_c_873_n 0.0101844f $X=5.54 $Y=2.815 $X2=0
+ $Y2=0
cc_516 N_A_515_392#_c_795_n N_VPWR_c_874_n 0.0129995f $X=6.44 $Y=2.455 $X2=0
+ $Y2=0
cc_517 N_A_515_392#_c_817_n N_VPWR_c_869_n 0.0093313f $X=5.425 $Y=2.385 $X2=0
+ $Y2=0
cc_518 N_A_515_392#_c_792_n N_VPWR_c_869_n 0.00842501f $X=5.54 $Y=2.815 $X2=0
+ $Y2=0
cc_519 N_A_515_392#_c_821_n N_VPWR_c_869_n 0.00923561f $X=6.275 $Y=2.385 $X2=0
+ $Y2=0
cc_520 N_A_515_392#_c_794_n N_VPWR_c_869_n 0.0100071f $X=4.61 $Y=2.465 $X2=0
+ $Y2=0
cc_521 N_A_515_392#_c_795_n N_VPWR_c_869_n 0.0121559f $X=6.44 $Y=2.455 $X2=0
+ $Y2=0
cc_522 N_VGND_c_941_n N_A_137_74#_c_1029_n 0.0111115f $X=0.295 $Y=0.49 $X2=0
+ $Y2=0
cc_523 N_VGND_c_942_n N_A_137_74#_c_1029_n 0.0106879f $X=2.115 $Y=0.515 $X2=0
+ $Y2=0
cc_524 N_VGND_c_944_n N_A_137_74#_c_1029_n 0.0460738f $X=1.95 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_948_n N_A_137_74#_c_1029_n 0.0386873f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_M1015_d N_A_593_74#_c_1044_n 0.00883733f $X=3.395 $Y=0.37 $X2=0
+ $Y2=0
cc_527 N_VGND_c_945_n N_A_593_74#_c_1044_n 0.0029521f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_c_946_n N_A_593_74#_c_1044_n 0.0029521f $X=5.385 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_c_948_n N_A_593_74#_c_1044_n 0.0115024f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_530 N_VGND_c_950_n N_A_593_74#_c_1044_n 0.0288883f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_531 N_VGND_c_945_n N_A_593_74#_c_1042_n 0.0105866f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_948_n N_A_593_74#_c_1042_n 0.00888607f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_c_950_n N_A_593_74#_c_1042_n 0.00283955f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_534 N_VGND_c_946_n N_A_593_74#_c_1043_n 0.0105866f $X=5.385 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_c_948_n N_A_593_74#_c_1043_n 0.00888607f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_950_n N_A_593_74#_c_1043_n 0.00283955f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_943_n N_A_981_74#_c_1068_n 0.0101711f $X=5.55 $Y=0.515 $X2=0
+ $Y2=0
cc_538 N_VGND_c_946_n N_A_981_74#_c_1068_n 0.0144296f $X=5.385 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_c_948_n N_A_981_74#_c_1068_n 0.0119645f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_540 N_VGND_M1000_d N_A_981_74#_c_1075_n 0.00353971f $X=5.405 $Y=0.37 $X2=0
+ $Y2=0
cc_541 N_VGND_c_943_n N_A_981_74#_c_1075_n 0.0166493f $X=5.55 $Y=0.515 $X2=0
+ $Y2=0
cc_542 N_VGND_c_948_n N_A_981_74#_c_1075_n 0.0123108f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_943_n N_A_981_74#_c_1069_n 0.0109329f $X=5.55 $Y=0.515 $X2=0
+ $Y2=0
cc_544 N_VGND_c_947_n N_A_981_74#_c_1069_n 0.0118609f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_c_948_n N_A_981_74#_c_1069_n 0.00912082f $X=6.48 $Y=0 $X2=0 $Y2=0
