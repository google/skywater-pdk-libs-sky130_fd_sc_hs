# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a2111oi_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a2111oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.450000 1.350000 8.035000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.205000 1.350000 9.555000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.350000 6.075000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 1.350000 3.510000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 1.180000 1.905000 1.550000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.708000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.840000 2.640000 1.010000 ;
        RECT 0.125000 1.010000 0.355000 1.720000 ;
        RECT 0.125000 1.720000 1.705000 1.890000 ;
        RECT 0.555000 1.890000 0.885000 2.735000 ;
        RECT 1.455000 1.890000 1.705000 2.735000 ;
        RECT 1.530000 0.330000 1.700000 0.840000 ;
        RECT 2.390000 0.350000 2.640000 0.840000 ;
        RECT 2.390000 1.010000 7.740000 1.130000 ;
        RECT 2.390000 1.130000 6.880000 1.180000 ;
        RECT 4.070000 0.350000 4.320000 0.975000 ;
        RECT 4.070000 0.975000 7.740000 1.010000 ;
        RECT 6.550000 0.770000 6.880000 0.915000 ;
        RECT 6.550000 0.915000 7.740000 0.975000 ;
        RECT 7.410000 0.770000 7.740000 0.915000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.105000  2.060000  0.355000 2.905000 ;
      RECT 0.105000  2.905000  2.235000 3.075000 ;
      RECT 1.020000  0.085000  1.350000 0.670000 ;
      RECT 1.085000  2.060000  1.255000 2.905000 ;
      RECT 1.880000  0.085000  2.210000 0.670000 ;
      RECT 1.905000  1.950000  4.035000 2.120000 ;
      RECT 1.905000  2.120000  2.235000 2.905000 ;
      RECT 2.435000  2.290000  2.685000 2.905000 ;
      RECT 2.435000  2.905000  5.925000 3.075000 ;
      RECT 2.810000  0.085000  3.900000 0.840000 ;
      RECT 2.855000  2.120000  3.085000 2.735000 ;
      RECT 3.255000  2.290000  3.585000 2.905000 ;
      RECT 3.705000  1.820000  4.035000 1.950000 ;
      RECT 3.755000  2.120000  4.035000 2.735000 ;
      RECT 4.245000  1.950000  9.975000 2.120000 ;
      RECT 4.245000  2.120000  4.525000 2.735000 ;
      RECT 4.500000  0.085000  4.830000 0.805000 ;
      RECT 4.695000  2.290000  5.025000 2.905000 ;
      RECT 5.195000  2.120000  5.425000 2.735000 ;
      RECT 5.595000  2.290000  5.925000 2.905000 ;
      RECT 6.120000  0.350000  8.090000 0.600000 ;
      RECT 6.120000  0.600000  6.380000 0.680000 ;
      RECT 6.125000  2.120000  6.295000 2.980000 ;
      RECT 6.495000  2.290000  6.825000 3.245000 ;
      RECT 7.025000  2.120000  7.195000 2.980000 ;
      RECT 7.040000  0.600000  7.250000 0.680000 ;
      RECT 7.395000  2.290000  7.725000 3.245000 ;
      RECT 7.920000  0.600000  8.090000 1.010000 ;
      RECT 7.920000  1.010000  9.890000 1.180000 ;
      RECT 7.925000  2.120000  8.095000 2.980000 ;
      RECT 8.270000  0.085000  8.600000 0.840000 ;
      RECT 8.295000  2.290000  8.545000 3.245000 ;
      RECT 8.745000  2.120000  9.075000 2.980000 ;
      RECT 8.780000  0.350000  8.950000 1.010000 ;
      RECT 9.130000  0.085000  9.460000 0.840000 ;
      RECT 9.275000  2.290000  9.525000 3.245000 ;
      RECT 9.640000  0.350000  9.890000 1.010000 ;
      RECT 9.725000  1.820000  9.975000 1.950000 ;
      RECT 9.725000  2.120000  9.975000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__a2111oi_4
END LIBRARY
