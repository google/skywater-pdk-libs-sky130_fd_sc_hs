* File: sky130_fd_sc_hs__o21a_2.spice
* Created: Tue Sep  1 20:14:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o21a_2.pex.spice"
.subckt sky130_fd_sc_hs__o21a_2  VNB VPB A1 A2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A1_M1006_g N_A_54_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1702 AS=0.2627 PD=1.2 PS=2.19 NRD=12.156 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1002 N_A_54_74#_M1002_d N_A2_M1002_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.1702 PD=1.065 PS=1.2 NRD=7.296 NRS=17.016 M=1 R=4.93333
+ SA=75000.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1009 N_A_244_368#_M1009_d N_B1_M1009_g N_A_54_74#_M1002_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.12025 PD=2.19 PS=1.065 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.4 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_X_M1000_d N_A_244_368#_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1000_d N_A_244_368#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 A_160_368# N_A1_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1004 N_A_244_368#_M1004_d N_A2_M1004_g A_160_368# VPB PSHORT L=0.15 W=1
+ AD=0.21 AS=0.135 PD=1.42 PS=1.27 NRD=25.5903 NRS=15.7403 M=1 R=6.66667
+ SA=75000.6 SB=75002 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_A_244_368#_M1004_d VPB PSHORT L=0.15 W=1
+ AD=0.276509 AS=0.21 PD=1.56604 PS=1.42 NRD=39.7152 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_244_368#_M1005_g N_VPWR_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.309691 PD=1.42 PS=1.75396 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1007 N_X_M1005_d N_A_244_368#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.2 SB=75000.3 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__o21a_2.pxi.spice"
*
.ends
*
*
