* File: sky130_fd_sc_hs__dlygate4sd3_1.spice
* Created: Tue Sep  1 20:03:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlygate4sd3_1.pex.spice"
.subckt sky130_fd_sc_hs__dlygate4sd3_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_28_74#_M1004_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1491 AS=0.1113 PD=1.13 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_A_289_74#_M1000_d N_A_28_74#_M1000_g N_VGND_M1004_d VNB NLOWVT L=0.18
+ W=0.42 AD=0.1092 AS=0.1491 PD=1.36 PS=1.13 NRD=0 NRS=107.136 M=1 R=2.33333
+ SA=90001 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1005 N_VGND_M1005_d N_A_289_74#_M1005_g N_A_405_138#_M1005_s VNB NLOWVT L=0.18
+ W=0.42 AD=0.0831672 AS=0.2436 PD=0.78569 PS=2 NRD=40.86 NRS=37.14 M=1
+ R=2.33333 SA=90000.5 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1006 N_X_M1006_d N_A_405_138#_M1006_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.146533 PD=2.01 PS=1.38431 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_28_74#_M1007_s VPB PSHORT L=0.15 W=0.42
+ AD=0.0894718 AS=0.1176 PD=0.81338 PS=1.4 NRD=14.0658 NRS=7.0329 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_A_289_74#_M1003_d N_A_28_74#_M1003_g N_VPWR_M1007_d VPB PSHORT L=0.5
+ W=1 AD=0.26 AS=0.213028 PD=2.52 PS=1.93662 NRD=0 NRS=12.7853 M=1 R=2 SA=250000
+ SB=250000 A=0.5 P=3 MULT=1
MM1001 N_VPWR_M1001_d N_A_289_74#_M1001_g N_A_405_138#_M1001_s VPB PSHORT L=0.5
+ W=1 AD=0.183019 AS=0.26 PD=1.39151 PS=2.52 NRD=13.2778 NRS=0 M=1 R=2 SA=250000
+ SB=250001 A=0.5 P=3 MULT=1
MM1002 N_X_M1002_d N_A_405_138#_M1002_g N_VPWR_M1001_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3136 AS=0.204981 PD=2.8 PS=1.55849 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__dlygate4sd3_1.pxi.spice"
*
.ends
*
*
