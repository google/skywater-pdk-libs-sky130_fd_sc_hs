* NGSPICE file created from sky130_fd_sc_hs__nand4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4_2 A B C D VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=2.268e+12p pd=1.525e+07u as=1.4112e+12p ps=1.148e+07u
M1001 a_515_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=6.2875e+11p pd=6.24e+06u as=2.22e+11p ps=2.08e+06u
M1002 Y B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y C VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR B Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=6.5035e+11p pd=6.28e+06u as=2.738e+11p ps=2.22e+06u
M1006 VPWR C Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y D VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_515_74# B a_304_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1009 a_304_74# C a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR D Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A a_515_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# C a_304_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_304_74# B a_515_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

