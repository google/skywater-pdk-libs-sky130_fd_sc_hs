* File: sky130_fd_sc_hs__sdfrtn_1.pex.spice
* Created: Tue Sep  1 20:22:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%SCE 3 6 7 9 12 15 22 23 25 26 27 33 35
c68 22 0 8.65763e-20 $X=0.7 $Y=1.575
r69 32 35 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.385 $Y=1.12
+ $X2=2.615 $Y2=1.12
r70 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.12 $X2=2.385 $Y2=1.12
r71 27 33 5.91467 $w=4.53e-07 $l=2.25e-07 $layer=LI1_cond $X=2.16 $Y=1.182
+ $X2=2.385 $Y2=1.182
r72 26 27 3.02306 $w=4.53e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=1.182
+ $X2=2.16 $Y2=1.182
r73 25 26 9.38335 $w=4.53e-07 $l=1.7e-07 $layer=LI1_cond $X=1.875 $Y=1.267
+ $X2=2.045 $Y2=1.267
r74 23 30 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.642 $Y=1.575
+ $X2=0.642 $Y2=1.41
r75 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.7
+ $Y=1.575 $X2=0.7 $Y2=1.575
r76 20 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=1.495
+ $X2=0.7 $Y2=1.495
r77 20 25 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.865 $Y=1.495
+ $X2=1.875 $Y2=1.495
r78 13 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=0.955
+ $X2=2.615 $Y2=1.12
r79 13 15 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.615 $Y=0.955
+ $X2=2.615 $Y2=0.615
r80 7 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.955 $Y=2.245
+ $X2=0.955 $Y2=2.64
r81 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r82 6 7 31.2407 $w=4.86e-07 $l=4.4477e-07 $layer=POLY_cond $X=0.642 $Y=1.93
+ $X2=0.955 $Y2=2.245
r83 5 23 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=0.642 $Y=1.632
+ $X2=0.642 $Y2=1.575
r84 5 6 37.2436 $w=4.45e-07 $l=2.98e-07 $layer=POLY_cond $X=0.642 $Y=1.632
+ $X2=0.642 $Y2=1.93
r85 3 30 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=0.65
+ $X2=0.495 $Y2=1.41
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_27_88# 1 2 9 11 12 14 17 20 23 25 31 32
+ 34 35 37 38 39 42
c92 11 0 1.86156e-19 $X=2.28 $Y=2.155
r93 38 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.1
+ $X2=1.455 $Y2=0.935
r94 37 39 7.86356 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=1.087
+ $X2=1.29 $Y2=1.087
r95 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.455
+ $Y=1.1 $X2=1.455 $Y2=1.1
r96 32 44 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.38 $Y=1.72 $X2=2.28
+ $Y2=1.72
r97 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.72 $X2=2.38 $Y2=1.72
r98 29 31 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=2.38 $Y=2.29
+ $X2=2.38 $Y2=1.72
r99 28 34 2.90107 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.145
+ $X2=0.28 $Y2=1.145
r100 28 39 49.3254 $w=1.88e-07 $l=8.45e-07 $layer=LI1_cond $X=0.445 $Y=1.145
+ $X2=1.29 $Y2=1.145
r101 26 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.375
+ $X2=0.24 $Y2=2.375
r102 25 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.215 $Y=2.375
+ $X2=2.38 $Y2=2.29
r103 25 26 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=2.215 $Y=2.375
+ $X2=0.365 $Y2=2.375
r104 21 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.375
r105 21 23 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.465
r106 20 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.29
+ $X2=0.24 $Y2=2.375
r107 19 34 3.58697 $w=2.9e-07 $l=1.13248e-07 $layer=LI1_cond $X=0.24 $Y=1.24
+ $X2=0.28 $Y2=1.145
r108 19 20 48.4026 $w=2.48e-07 $l=1.05e-06 $layer=LI1_cond $X=0.24 $Y=1.24
+ $X2=0.24 $Y2=2.29
r109 15 34 3.58697 $w=2.9e-07 $l=9.5e-08 $layer=LI1_cond $X=0.28 $Y=1.05
+ $X2=0.28 $Y2=1.145
r110 15 17 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.28 $Y=1.05 $X2=0.28
+ $Y2=0.65
r111 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.28 $Y=2.245
+ $X2=2.28 $Y2=2.64
r112 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.28 $Y=2.155
+ $X2=2.28 $Y2=2.245
r113 10 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.885
+ $X2=2.28 $Y2=1.72
r114 10 11 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.28 $Y=1.885
+ $X2=2.28 $Y2=2.155
r115 9 42 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.545 $Y=0.615
+ $X2=1.545 $Y2=0.935
r116 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r117 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.44 $X2=0.28 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%D 1 3 4 8 10 12 13 17 18
c40 18 0 1.86156e-19 $X=1.815 $Y=1.945
c41 10 0 8.65763e-20 $X=1.345 $Y=2.035
r42 17 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.815 $Y=1.945
+ $X2=1.815 $Y2=2.035
r43 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.945
+ $X2=1.815 $Y2=1.78
r44 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.815
+ $Y=1.945 $X2=1.815 $Y2=1.945
r45 13 18 4.57588 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.68 $Y=1.95
+ $X2=1.815 $Y2=1.95
r46 12 13 16.2698 $w=3.38e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.95 $X2=1.68
+ $Y2=1.95
r47 8 19 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=1.905 $Y=0.615
+ $X2=1.905 $Y2=1.78
r48 5 10 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.435 $Y=2.035 $X2=1.345
+ $Y2=2.035
r49 4 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=2.035
+ $X2=1.815 $Y2=2.035
r50 4 5 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.65 $Y=2.035
+ $X2=1.435 $Y2=2.035
r51 1 10 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=1.345 $Y=2.245
+ $X2=1.345 $Y2=2.035
r52 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.345 $Y=2.245
+ $X2=1.345 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%SCD 1 3 5 8 12 14 15 19
c50 5 0 1.38402e-19 $X=2.875 $Y=2.095
r51 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.69
+ $X2=2.965 $Y2=1.855
r52 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.69
+ $X2=2.965 $Y2=1.525
r53 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.69 $X2=2.965 $Y2=1.69
r54 15 20 9.14007 $w=4.33e-07 $l=3.45e-07 $layer=LI1_cond $X=3.017 $Y=2.035
+ $X2=3.017 $Y2=1.69
r55 14 20 0.662324 $w=4.33e-07 $l=2.5e-08 $layer=LI1_cond $X=3.017 $Y=1.665
+ $X2=3.017 $Y2=1.69
r56 10 12 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.67 $Y=2.17
+ $X2=2.875 $Y2=2.17
r57 8 21 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.005 $Y=0.615
+ $X2=3.005 $Y2=1.525
r58 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=2.095
+ $X2=2.875 $Y2=2.17
r59 5 22 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.875 $Y=2.095
+ $X2=2.875 $Y2=1.855
r60 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=2.245
+ $X2=2.67 $Y2=2.17
r61 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.67 $Y=2.245
+ $X2=2.67 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%RESET_B 1 3 6 9 10 12 15 18 21 24 25 27 28
+ 30 31 32 33 38 41 44 45 48 49 53 54
c216 53 0 1.97052e-19 $X=11.16 $Y=1.375
c217 49 0 8.36181e-20 $X=7.85 $Y=1.635
c218 48 0 1.0834e-19 $X=7.85 $Y=1.635
c219 45 0 1.38402e-19 $X=3.57 $Y=1.52
c220 30 0 1.8853e-19 $X=7.775 $Y=1.665
c221 28 0 2.78046e-19 $X=11.25 $Y=2.375
r222 53 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.16 $Y=1.375
+ $X2=11.16 $Y2=1.54
r223 53 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.16 $Y=1.375
+ $X2=11.16 $Y2=1.21
r224 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.16
+ $Y=1.375 $X2=11.16 $Y2=1.375
r225 48 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.85 $Y=1.635
+ $X2=7.85 $Y2=1.8
r226 48 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.85 $Y=1.635
+ $X2=7.85 $Y2=1.47
r227 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.85
+ $Y=1.635 $X2=7.85 $Y2=1.635
r228 44 46 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.552 $Y=1.52
+ $X2=3.552 $Y2=1.355
r229 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.52 $X2=3.57 $Y2=1.52
r230 41 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=1.665
+ $X2=3.6 $Y2=1.665
r231 39 54 11.2317 $w=3.15e-07 $l=2.9e-07 $layer=LI1_cond $X=11.195 $Y=1.665
+ $X2=11.195 $Y2=1.375
r232 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=1.665
+ $X2=11.28 $Y2=1.665
r233 35 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.665
r234 33 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=1.665
+ $X2=7.92 $Y2=1.665
r235 32 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.135 $Y=1.665
+ $X2=11.28 $Y2=1.665
r236 32 33 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=11.135 $Y=1.665
+ $X2=8.065 $Y2=1.665
r237 31 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=1.665
+ $X2=3.6 $Y2=1.665
r238 30 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=1.665
+ $X2=7.92 $Y2=1.665
r239 30 31 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=7.775 $Y=1.665
+ $X2=3.745 $Y2=1.665
r240 28 29 19.6163 $w=1.72e-07 $l=7e-08 $layer=POLY_cond $X=11.25 $Y=2.375
+ $X2=11.32 $Y2=2.375
r241 25 29 6.07713 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.32 $Y=2.465
+ $X2=11.32 $Y2=2.375
r242 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.32 $Y=2.465
+ $X2=11.32 $Y2=2.75
r243 24 28 6.07713 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.25 $Y=2.285
+ $X2=11.25 $Y2=2.375
r244 24 56 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=11.25 $Y=2.285
+ $X2=11.25 $Y2=1.54
r245 21 55 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=11.25 $Y=0.58
+ $X2=11.25 $Y2=1.21
r246 18 51 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.79 $Y=2.11
+ $X2=7.79 $Y2=1.8
r247 15 50 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=7.76 $Y=0.865
+ $X2=7.76 $Y2=1.47
r248 10 18 78.4908 $w=2.18e-07 $l=4.04104e-07 $layer=POLY_cond $X=7.685 $Y=2.465
+ $X2=7.79 $Y2=2.11
r249 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.685 $Y=2.465
+ $X2=7.685 $Y2=2.75
r250 8 44 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=3.552 $Y=1.537
+ $X2=3.552 $Y2=1.52
r251 8 9 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=3.552 $Y=1.537
+ $X2=3.552 $Y2=1.843
r252 6 46 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.445 $Y=0.615
+ $X2=3.445 $Y2=1.355
r253 1 9 62.5045 $w=3.1e-07 $l=5.16651e-07 $layer=POLY_cond $X=3.29 $Y=2.245
+ $X2=3.552 $Y2=1.843
r254 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.29 $Y=2.245
+ $X2=3.29 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%CLK_N 1 3 4 6 7
c37 4 0 1.90908e-19 $X=4.375 $Y=1.765
r38 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.44
+ $Y=1.385 $X2=4.44 $Y2=1.385
r39 7 11 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=4.56 $Y=1.38 $X2=4.44
+ $Y2=1.38
r40 4 10 67.4361 $w=3.64e-07 $l=3.86445e-07 $layer=POLY_cond $X=4.375 $Y=1.765
+ $X2=4.362 $Y2=1.385
r41 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.375 $Y=1.765
+ $X2=4.375 $Y2=2.4
r42 1 10 38.9663 $w=3.64e-07 $l=2.35465e-07 $layer=POLY_cond $X=4.195 $Y=1.22
+ $X2=4.362 $Y2=1.385
r43 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.195 $Y=1.22 $X2=4.195
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_1074_88# 1 2 7 9 11 12 14 16 17 19 20 22
+ 24 25 28 31 32 36 37 38 41 42 43 44 48 50 54 55 67
c183 50 0 9.45937e-20 $X=6.26 $Y=1.94
c184 48 0 1.72856e-19 $X=6.425 $Y=1.94
c185 25 0 1.14899e-19 $X=6.755 $Y=1.94
c186 11 0 1.32863e-19 $X=6.845 $Y=2.375
r187 59 70 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.66 $Y=1.065
+ $X2=9.66 $Y2=1.23
r188 59 67 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=9.66 $Y=1.065
+ $X2=9.66 $Y2=0.94
r189 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.66
+ $Y=1.065 $X2=9.66 $Y2=1.065
r190 55 58 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.66 $Y=0.875
+ $X2=9.66 $Y2=1.065
r191 54 63 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.49 $Y=0.38
+ $X2=6.285 $Y2=0.38
r192 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.49
+ $Y=0.38 $X2=6.49 $Y2=0.38
r193 48 50 6.00814 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=1.94
+ $X2=6.26 $Y2=1.94
r194 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.425
+ $Y=1.94 $X2=6.425 $Y2=1.94
r195 42 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=0.875
+ $X2=9.66 $Y2=0.875
r196 42 43 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=9.495 $Y=0.875
+ $X2=7.27 $Y2=0.875
r197 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.185 $Y=0.79
+ $X2=7.27 $Y2=0.875
r198 40 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.185 $Y=0.545
+ $X2=7.185 $Y2=0.79
r199 39 53 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.495 $Y=0.4
+ $X2=6.41 $Y2=0.4
r200 38 40 7.43784 $w=2.9e-07 $l=1.8262e-07 $layer=LI1_cond $X=7.1 $Y=0.4
+ $X2=7.185 $Y2=0.545
r201 38 39 24.0423 $w=2.88e-07 $l=6.05e-07 $layer=LI1_cond $X=7.1 $Y=0.4
+ $X2=6.495 $Y2=0.4
r202 36 53 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.41 $Y=0.545
+ $X2=6.41 $Y2=0.4
r203 36 37 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.41 $Y=0.545
+ $X2=6.41 $Y2=1.265
r204 35 46 3.61267 $w=2.85e-07 $l=2.22374e-07 $layer=LI1_cond $X=5.775 $Y=1.962
+ $X2=5.56 $Y2=1.977
r205 35 50 19.6117 $w=2.83e-07 $l=4.85e-07 $layer=LI1_cond $X=5.775 $Y=1.962
+ $X2=6.26 $Y2=1.962
r206 33 44 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.675 $Y=1.35
+ $X2=5.51 $Y2=1.35
r207 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.325 $Y=1.35
+ $X2=6.41 $Y2=1.265
r208 32 33 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.325 $Y=1.35
+ $X2=5.675 $Y2=1.35
r209 31 46 3.2514 $w=3.3e-07 $l=1.80275e-07 $layer=LI1_cond $X=5.51 $Y=1.82
+ $X2=5.56 $Y2=1.977
r210 30 44 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.51 $Y=1.435
+ $X2=5.51 $Y2=1.35
r211 30 31 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.51 $Y=1.435
+ $X2=5.51 $Y2=1.82
r212 26 44 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.51 $Y=1.265
+ $X2=5.51 $Y2=1.35
r213 26 28 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.51 $Y=1.265
+ $X2=5.51 $Y2=1.035
r214 25 49 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=6.755 $Y=1.94
+ $X2=6.425 $Y2=1.94
r215 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.29 $Y=0.865
+ $X2=10.29 $Y2=0.58
r216 21 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.825 $Y=0.94
+ $X2=9.66 $Y2=0.94
r217 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.215 $Y=0.94
+ $X2=10.29 $Y2=0.865
r218 20 21 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=10.215 $Y=0.94
+ $X2=9.825 $Y2=0.94
r219 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.62 $Y=1.885
+ $X2=9.62 $Y2=2.46
r220 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.62 $Y=1.795
+ $X2=9.62 $Y2=1.885
r221 16 70 219.621 $w=1.8e-07 $l=5.65e-07 $layer=POLY_cond $X=9.62 $Y=1.795
+ $X2=9.62 $Y2=1.23
r222 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.845 $Y=2.465
+ $X2=6.845 $Y2=2.75
r223 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.845 $Y=2.375
+ $X2=6.845 $Y2=2.465
r224 10 25 14.8326 $w=5.17e-07 $l=2.96606e-07 $layer=POLY_cond $X=6.845 $Y=2.195
+ $X2=6.755 $Y2=1.94
r225 10 11 69.9677 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=6.845 $Y=2.195
+ $X2=6.845 $Y2=2.375
r226 7 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.285 $Y=0.545
+ $X2=6.285 $Y2=0.38
r227 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.285 $Y=0.545
+ $X2=6.285 $Y2=0.865
r228 2 46 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.84 $X2=5.61 $Y2=2.015
r229 1 28 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.37
+ $Y=0.44 $X2=5.51 $Y2=1.035
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_1429_308# 1 2 8 9 11 14 18 19 21 22 23 27
+ 32 33
c98 32 0 1.69146e-19 $X=8.96 $Y=2.135
c99 18 0 1.14899e-19 $X=7.31 $Y=1.705
c100 14 0 8.36181e-20 $X=7.37 $Y=0.865
r101 32 34 0.276272 $w=8.73e-07 $l=5e-09 $layer=LI1_cond $X=9.127 $Y=2.135
+ $X2=9.127 $Y2=2.14
r102 32 33 12.1237 $w=8.73e-07 $l=1.65e-07 $layer=LI1_cond $X=9.127 $Y=2.135
+ $X2=9.127 $Y2=1.97
r103 27 34 10.4851 $w=7.68e-07 $l=6.75e-07 $layer=LI1_cond $X=9.18 $Y=2.815
+ $X2=9.18 $Y2=2.14
r104 23 30 3.40825 $w=1.7e-07 $l=1.16619e-07 $layer=LI1_cond $X=8.775 $Y=1.3
+ $X2=8.85 $Y2=1.215
r105 23 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.775 $Y=1.3
+ $X2=8.775 $Y2=1.97
r106 21 30 3.40825 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.69 $Y=1.215
+ $X2=8.85 $Y2=1.215
r107 21 22 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=8.69 $Y=1.215
+ $X2=7.475 $Y2=1.215
r108 19 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.31 $Y=1.705
+ $X2=7.31 $Y2=1.87
r109 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.31 $Y=1.705
+ $X2=7.31 $Y2=1.54
r110 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.705 $X2=7.31 $Y2=1.705
r111 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.31 $Y=1.3
+ $X2=7.475 $Y2=1.215
r112 16 18 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=7.31 $Y=1.3
+ $X2=7.31 $Y2=1.705
r113 14 36 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=7.37 $Y=0.865
+ $X2=7.37 $Y2=1.54
r114 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.235 $Y=2.465
+ $X2=7.235 $Y2=2.75
r115 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.235 $Y=2.375
+ $X2=7.235 $Y2=2.465
r116 8 37 196.298 $w=1.8e-07 $l=5.05e-07 $layer=POLY_cond $X=7.235 $Y=2.375
+ $X2=7.235 $Y2=1.87
r117 2 32 200 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=3 $X=8.76
+ $Y=1.96 $X2=8.96 $Y2=2.135
r118 2 27 200 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=3 $X=8.76
+ $Y=1.96 $X2=8.96 $Y2=2.815
r119 1 30 182 $w=1.7e-07 $l=6.19375e-07 $layer=licon1_NDIFF $count=1 $X=8.425
+ $Y=0.72 $X2=8.705 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_1272_131# 1 2 3 10 12 13 15 18 21 22 24
+ 26 30 31 33 37
c111 30 0 7.49297e-20 $X=8.39 $Y=1.635
c112 24 0 1.8853e-19 $X=7.91 $Y=2.445
c113 22 0 1.0834e-19 $X=7.745 $Y=2.36
r114 35 37 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.755 $Y=0.93
+ $X2=6.845 $Y2=0.93
r115 31 43 39.8291 $w=3.57e-07 $l=2.95e-07 $layer=POLY_cond $X=8.39 $Y=1.677
+ $X2=8.685 $Y2=1.677
r116 31 41 5.40056 $w=3.57e-07 $l=4e-08 $layer=POLY_cond $X=8.39 $Y=1.677
+ $X2=8.35 $Y2=1.677
r117 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.39
+ $Y=1.635 $X2=8.39 $Y2=1.635
r118 28 30 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=8.372 $Y=1.97
+ $X2=8.372 $Y2=1.635
r119 24 28 23.8831 $w=2.36e-07 $l=6.01837e-07 $layer=LI1_cond $X=7.91 $Y=2.292
+ $X2=8.372 $Y2=1.97
r120 24 26 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=7.91 $Y=2.445
+ $X2=7.91 $Y2=2.75
r121 23 33 2.76166 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=6.93 $Y=2.36
+ $X2=6.692 $Y2=2.36
r122 22 24 9.50365 $w=2.36e-07 $l=1.96074e-07 $layer=LI1_cond $X=7.745 $Y=2.36
+ $X2=7.91 $Y2=2.292
r123 22 23 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=7.745 $Y=2.36
+ $X2=6.93 $Y2=2.36
r124 21 33 3.70735 $w=2.5e-07 $l=1.90825e-07 $layer=LI1_cond $X=6.845 $Y=2.275
+ $X2=6.692 $Y2=2.36
r125 20 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=1.095
+ $X2=6.845 $Y2=0.93
r126 20 21 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=6.845 $Y=1.095
+ $X2=6.845 $Y2=2.275
r127 16 33 3.70735 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=6.62 $Y=2.445
+ $X2=6.692 $Y2=2.36
r128 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.62 $Y=2.445
+ $X2=6.62 $Y2=2.75
r129 13 43 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.685 $Y=1.885
+ $X2=8.685 $Y2=1.677
r130 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.685 $Y=1.885
+ $X2=8.685 $Y2=2.46
r131 10 41 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.35 $Y=1.47
+ $X2=8.35 $Y2=1.677
r132 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.35 $Y=1.47
+ $X2=8.35 $Y2=1.04
r133 3 26 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.54 $X2=7.91 $Y2=2.75
r134 2 18 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=6.47
+ $Y=2.54 $X2=6.62 $Y2=2.75
r135 1 35 182 $w=1.7e-07 $l=5.14441e-07 $layer=licon1_NDIFF $count=1 $X=6.36
+ $Y=0.655 $X2=6.755 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_854_74# 1 2 7 9 10 12 13 14 16 17 19 20
+ 21 23 24 29 30 31 35 37 38 40 41 44 45 49 53 60 64 66 68 71 73 74 75
c213 37 0 1.69146e-19 $X=10.135 $Y=2.375
c214 16 0 1.72856e-19 $X=5.945 $Y=2.315
c215 13 0 9.45937e-20 $X=5.87 $Y=1.49
r216 74 83 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=10.23 $Y=1.39
+ $X2=10.135 $Y2=1.39
r217 73 75 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=10.23 $Y=1.382
+ $X2=10.065 $Y2=1.382
r218 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.23
+ $Y=1.39 $X2=10.23 $Y2=1.39
r219 71 79 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=9.155 $Y=1.635
+ $X2=9.06 $Y2=1.635
r220 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.155
+ $Y=1.635 $X2=9.155 $Y2=1.635
r221 68 70 7.70526 $w=2.85e-07 $l=1.8e-07 $layer=LI1_cond $X=9.19 $Y=1.455
+ $X2=9.19 $Y2=1.635
r222 64 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.01 $Y=1.455
+ $X2=5.01 $Y2=1.62
r223 64 66 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.01 $Y=1.455
+ $X2=5.01 $Y2=1.29
r224 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=1.455 $X2=5.01 $Y2=1.455
r225 62 68 3.76007 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=9.35 $Y=1.455
+ $X2=9.19 $Y2=1.455
r226 62 75 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.35 $Y=1.455
+ $X2=10.065 $Y2=1.455
r227 60 67 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.93 $Y=1.82 $X2=4.93
+ $Y2=1.62
r228 57 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.93 $Y=1.04
+ $X2=4.93 $Y2=1.29
r229 53 60 7.64049 $w=3.15e-07 $l=1.94921e-07 $layer=LI1_cond $X=4.845 $Y=1.977
+ $X2=4.93 $Y2=1.82
r230 53 55 8.96345 $w=3.13e-07 $l=2.45e-07 $layer=LI1_cond $X=4.845 $Y=1.977
+ $X2=4.6 $Y2=1.977
r231 49 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.845 $Y=0.955
+ $X2=4.93 $Y2=1.04
r232 49 51 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.845 $Y=0.955
+ $X2=4.41 $Y2=0.955
r233 45 47 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=6.675 $Y=1.225
+ $X2=6.675 $Y2=1.49
r234 42 43 10.0417 $w=4.32e-07 $l=9e-08 $layer=POLY_cond $X=5.295 $Y=1.527
+ $X2=5.385 $Y2=1.527
r235 41 65 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.22 $Y=1.455
+ $X2=5.01 $Y2=1.455
r236 41 42 11.1745 $w=4.32e-07 $l=1.05e-07 $layer=POLY_cond $X=5.22 $Y=1.455
+ $X2=5.295 $Y2=1.527
r237 38 40 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.135 $Y=2.465
+ $X2=10.135 $Y2=2.75
r238 37 38 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.135 $Y=2.375
+ $X2=10.135 $Y2=2.465
r239 36 83 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.135 $Y=1.555
+ $X2=10.135 $Y2=1.39
r240 36 37 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=10.135 $Y=1.555
+ $X2=10.135 $Y2=2.375
r241 33 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.06 $Y=1.47
+ $X2=9.06 $Y2=1.635
r242 33 35 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.06 $Y=1.47
+ $X2=9.06 $Y2=1.04
r243 32 35 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=9.06 $Y=0.285
+ $X2=9.06 $Y2=1.04
r244 30 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.985 $Y=0.21
+ $X2=9.06 $Y2=0.285
r245 30 31 989.638 $w=1.5e-07 $l=1.93e-06 $layer=POLY_cond $X=8.985 $Y=0.21
+ $X2=7.055 $Y2=0.21
r246 27 29 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.98 $Y=1.15
+ $X2=6.98 $Y2=0.865
r247 26 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.98 $Y=0.285
+ $X2=7.055 $Y2=0.21
r248 26 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.98 $Y=0.285
+ $X2=6.98 $Y2=0.865
r249 25 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.75 $Y=1.225
+ $X2=6.675 $Y2=1.225
r250 24 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.905 $Y=1.225
+ $X2=6.98 $Y2=1.15
r251 24 25 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=6.905 $Y=1.225
+ $X2=6.75 $Y2=1.225
r252 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.395 $Y=2.465
+ $X2=6.395 $Y2=2.75
r253 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.32 $Y=2.39
+ $X2=6.395 $Y2=2.465
r254 19 20 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=6.32 $Y=2.39 $X2=6.02
+ $Y2=2.39
r255 18 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.02 $Y=1.49
+ $X2=5.945 $Y2=1.49
r256 17 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.6 $Y=1.49
+ $X2=6.675 $Y2=1.49
r257 17 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.6 $Y=1.49
+ $X2=6.02 $Y2=1.49
r258 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.945 $Y=2.315
+ $X2=6.02 $Y2=2.39
r259 15 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.945 $Y=1.565
+ $X2=5.945 $Y2=1.49
r260 15 16 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.945 $Y=1.565
+ $X2=5.945 $Y2=2.315
r261 14 43 31.8951 $w=4.32e-07 $l=1.06911e-07 $layer=POLY_cond $X=5.475 $Y=1.49
+ $X2=5.385 $Y2=1.527
r262 13 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.87 $Y=1.49
+ $X2=5.945 $Y2=1.49
r263 13 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.87 $Y=1.49
+ $X2=5.475 $Y2=1.49
r264 10 43 27.7542 $w=1.5e-07 $l=2.38e-07 $layer=POLY_cond $X=5.385 $Y=1.765
+ $X2=5.385 $Y2=1.527
r265 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.385 $Y=1.765
+ $X2=5.385 $Y2=2.4
r266 7 42 27.7542 $w=1.5e-07 $l=2.37e-07 $layer=POLY_cond $X=5.295 $Y=1.29
+ $X2=5.295 $Y2=1.527
r267 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.295 $Y=1.29
+ $X2=5.295 $Y2=0.81
r268 2 55 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=4.45
+ $Y=1.84 $X2=4.6 $Y2=2.015
r269 1 51 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.37 $X2=4.41 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_2087_410# 1 2 7 9 12 14 18 20 24 27 29 34
c91 29 0 9.65573e-20 $X=10.6 $Y=2.215
c92 12 0 1.91401e-20 $X=10.69 $Y=0.58
r93 29 32 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=10.56 $Y=2.215
+ $X2=10.56 $Y2=2.375
r94 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.6
+ $Y=2.215 $X2=10.6 $Y2=2.215
r95 26 27 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=12.15 $Y=0.7
+ $X2=12.15 $Y2=2.29
r96 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.71 $Y=2.375
+ $X2=11.545 $Y2=2.375
r97 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.065 $Y=2.375
+ $X2=12.15 $Y2=2.29
r98 24 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.065 $Y=2.375
+ $X2=11.71 $Y2=2.375
r99 20 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.065 $Y=0.575
+ $X2=12.15 $Y2=0.7
r100 20 22 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=12.065 $Y=0.575
+ $X2=11.96 $Y2=0.575
r101 16 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.545 $Y=2.46
+ $X2=11.545 $Y2=2.375
r102 16 18 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=11.545 $Y=2.46
+ $X2=11.545 $Y2=2.75
r103 15 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.685 $Y=2.375
+ $X2=10.56 $Y2=2.375
r104 14 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.38 $Y=2.375
+ $X2=11.545 $Y2=2.375
r105 14 15 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=11.38 $Y=2.375
+ $X2=10.685 $Y2=2.375
r106 10 30 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=10.69 $Y=2.05
+ $X2=10.6 $Y2=2.215
r107 10 12 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=10.69 $Y=2.05
+ $X2=10.69 $Y2=0.58
r108 7 30 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=10.545 $Y=2.465
+ $X2=10.6 $Y2=2.215
r109 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.545 $Y=2.465
+ $X2=10.545 $Y2=2.75
r110 2 18 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.395
+ $Y=2.54 $X2=11.545 $Y2=2.75
r111 1 22 182 $w=1.7e-07 $l=3.46482e-07 $layer=licon1_NDIFF $count=1 $X=11.715
+ $Y=0.37 $X2=11.96 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_1827_144# 1 2 7 9 11 13 15 16 18 19 21 23
+ 25 26 28 29 30 35 39 40 41 42 43 44 45 50 51 53 54
c159 54 0 1.97052e-19 $X=10.94 $Y=1.795
c160 40 0 1.91401e-20 $X=10.08 $Y=0.87
c161 21 0 1.07922e-19 $X=12.77 $Y=1.07
c162 19 0 1.07922e-19 $X=12.755 $Y=1.97
r163 54 56 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.94 $Y=1.795
+ $X2=10.94 $Y2=2.035
r164 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.73
+ $Y=1.065 $X2=11.73 $Y2=1.065
r165 48 50 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=11.73 $Y=1.95
+ $X2=11.73 $Y2=1.065
r166 47 50 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=11.73 $Y=1.04
+ $X2=11.73 $Y2=1.065
r167 46 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.025 $Y=2.035
+ $X2=10.94 $Y2=2.035
r168 45 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.565 $Y=2.035
+ $X2=11.73 $Y2=1.95
r169 45 46 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=11.565 $Y=2.035
+ $X2=11.025 $Y2=2.035
r170 43 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.565 $Y=0.955
+ $X2=11.73 $Y2=1.04
r171 43 44 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=11.565 $Y=0.955
+ $X2=10.165 $Y2=0.955
r172 41 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.855 $Y=1.795
+ $X2=10.94 $Y2=1.795
r173 41 42 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=10.855 $Y=1.795
+ $X2=10.065 $Y2=1.795
r174 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.08 $Y=0.87
+ $X2=10.165 $Y2=0.955
r175 39 53 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.08 $Y=0.62
+ $X2=10.08 $Y2=0.455
r176 39 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=10.08 $Y=0.62
+ $X2=10.08 $Y2=0.87
r177 35 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.9 $Y=2.135
+ $X2=9.9 $Y2=2.815
r178 33 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.9 $Y=1.88
+ $X2=10.065 $Y2=1.795
r179 33 35 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.9 $Y=1.88
+ $X2=9.9 $Y2=2.135
r180 26 28 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=12.845 $Y=0.995
+ $X2=12.845 $Y2=0.645
r181 23 25 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.83 $Y=2.045
+ $X2=12.83 $Y2=2.54
r182 22 51 12.1617 $w=1.5e-07 $l=1.8747e-07 $layer=POLY_cond $X=11.895 $Y=1.07
+ $X2=11.73 $Y2=1.022
r183 21 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.77 $Y=1.07
+ $X2=12.845 $Y2=0.995
r184 21 22 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=12.77 $Y=1.07
+ $X2=11.895 $Y2=1.07
r185 20 30 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.86 $Y=1.97
+ $X2=11.77 $Y2=1.97
r186 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.755 $Y=1.97
+ $X2=12.83 $Y2=2.045
r187 19 20 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=12.755 $Y=1.97
+ $X2=11.86 $Y2=1.97
r188 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.77 $Y=2.465
+ $X2=11.77 $Y2=2.75
r189 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.77 $Y=2.375
+ $X2=11.77 $Y2=2.465
r190 14 30 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.77 $Y=2.045
+ $X2=11.77 $Y2=1.97
r191 14 15 128.274 $w=1.8e-07 $l=3.3e-07 $layer=POLY_cond $X=11.77 $Y=2.045
+ $X2=11.77 $Y2=2.375
r192 13 30 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.755
+ $Y=1.895 $X2=11.77 $Y2=1.97
r193 13 29 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=11.755 $Y=1.895
+ $X2=11.755 $Y2=1.57
r194 11 29 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.73 $Y=1.405
+ $X2=11.73 $Y2=1.57
r195 10 51 13.5877 $w=2.4e-07 $l=1.23e-07 $layer=POLY_cond $X=11.73 $Y=1.145
+ $X2=11.73 $Y2=1.022
r196 10 11 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=11.73 $Y=1.145
+ $X2=11.73 $Y2=1.405
r197 7 51 13.5877 $w=2.4e-07 $l=1.60823e-07 $layer=POLY_cond $X=11.64 $Y=0.9
+ $X2=11.73 $Y2=1.022
r198 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.64 $Y=0.9
+ $X2=11.64 $Y2=0.58
r199 2 37 600 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=9.695
+ $Y=1.96 $X2=9.9 $Y2=2.815
r200 2 35 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=9.695
+ $Y=1.96 $X2=9.845 $Y2=2.135
r201 1 53 91 $w=1.7e-07 $l=9.83616e-07 $layer=licon1_NDIFF $count=2 $X=9.135
+ $Y=0.72 $X2=9.995 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_2492_424# 1 2 7 9 12 14 15 18 22 25
c45 25 0 2.15844e-19 $X=12.645 $Y=1.52
r46 25 28 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.625 $Y=1.52
+ $X2=12.625 $Y2=1.685
r47 25 27 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.625 $Y=1.52
+ $X2=12.625 $Y2=1.355
r48 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.645
+ $Y=1.52 $X2=12.645 $Y2=1.52
r49 22 28 18.8286 $w=3.53e-07 $l=5.8e-07 $layer=LI1_cond $X=12.617 $Y=2.265
+ $X2=12.617 $Y2=1.685
r50 18 27 23.0489 $w=3.53e-07 $l=7.1e-07 $layer=LI1_cond $X=12.617 $Y=0.645
+ $X2=12.617 $Y2=1.355
r51 14 26 118.031 $w=3.3e-07 $l=6.75e-07 $layer=POLY_cond $X=13.32 $Y=1.52
+ $X2=12.645 $Y2=1.52
r52 14 15 5.03009 $w=3.3e-07 $l=1.08167e-07 $layer=POLY_cond $X=13.32 $Y=1.52
+ $X2=13.41 $Y2=1.56
r53 10 15 37.0704 $w=1.5e-07 $l=2.12368e-07 $layer=POLY_cond $X=13.425 $Y=1.355
+ $X2=13.41 $Y2=1.56
r54 10 12 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=13.425 $Y=1.355
+ $X2=13.425 $Y2=0.74
r55 7 15 37.0704 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=13.41 $Y=1.765
+ $X2=13.41 $Y2=1.56
r56 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.41 $Y=1.765
+ $X2=13.41 $Y2=2.4
r57 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=12.46
+ $Y=2.12 $X2=12.605 $Y2=2.265
r58 1 18 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=12.485
+ $Y=0.37 $X2=12.63 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 36 40 44 48 52
+ 56 61 64 68 69 70 72 84 88 96 101 113 119 120 123 126 129 132 135 138 145
c156 138 0 1.81488e-19 $X=10.905 $Y=2.815
c157 6 0 7.49297e-20 $X=8.325 $Y=1.96
r158 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r159 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r160 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r161 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r162 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r163 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r164 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r165 120 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r166 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r167 117 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=3.33
+ $X2=13.14 $Y2=3.33
r168 117 119 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.305 $Y=3.33
+ $X2=13.68 $Y2=3.33
r169 116 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r170 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r171 113 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=3.33
+ $X2=13.14 $Y2=3.33
r172 113 115 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.975 $Y=3.33
+ $X2=12.72 $Y2=3.33
r173 112 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r174 112 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r175 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r176 109 111 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=11.21 $Y=3.33
+ $X2=11.76 $Y2=3.33
r177 108 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r178 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r179 105 108 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r180 105 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r181 104 107 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r182 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r183 102 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.46 $Y2=3.33
r184 102 104 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.88 $Y2=3.33
r185 101 109 8.37032 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=10.907 $Y=3.33
+ $X2=11.21 $Y2=3.33
r186 101 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r187 101 138 10.1815 $w=6.03e-07 $l=5.15e-07 $layer=LI1_cond $X=10.907 $Y=3.33
+ $X2=10.907 $Y2=2.815
r188 101 107 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.605 $Y=3.33
+ $X2=10.32 $Y2=3.33
r189 100 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r190 100 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r191 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r192 97 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.42 $Y2=3.33
r193 97 99 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.92 $Y2=3.33
r194 96 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.46 $Y2=3.33
r195 96 99 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=7.92 $Y2=3.33
r196 92 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r197 91 94 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.96 $Y2=3.33
r198 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r199 89 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=3.33
+ $X2=5.16 $Y2=3.33
r200 89 91 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.325 $Y=3.33
+ $X2=5.52 $Y2=3.33
r201 88 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.295 $Y=3.33
+ $X2=7.42 $Y2=3.33
r202 88 94 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.295 $Y=3.33
+ $X2=6.96 $Y2=3.33
r203 87 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r204 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r205 84 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=3.33
+ $X2=4.075 $Y2=3.33
r206 84 86 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.91 $Y=3.33
+ $X2=3.6 $Y2=3.33
r207 83 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r208 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r209 80 83 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r210 80 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r211 79 82 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r212 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r213 77 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r214 77 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r215 75 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r216 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r217 72 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r218 72 74 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r219 70 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r220 70 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=5.52 $Y2=3.33
r221 70 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r222 68 111 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=11.88 $Y=3.33
+ $X2=11.76 $Y2=3.33
r223 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.88 $Y=3.33
+ $X2=12.045 $Y2=3.33
r224 67 115 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=12.21 $Y=3.33
+ $X2=12.72 $Y2=3.33
r225 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.21 $Y=3.33
+ $X2=12.045 $Y2=3.33
r226 65 86 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=3.6 $Y2=3.33
r227 64 82 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.64 $Y2=3.33
r228 63 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.98 $Y=3.33
+ $X2=3.145 $Y2=3.33
r229 63 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.98 $Y=3.33
+ $X2=2.815 $Y2=3.33
r230 61 63 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.98 $Y=3.055
+ $X2=2.98 $Y2=3.33
r231 56 59 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=13.14 $Y=1.985
+ $X2=13.14 $Y2=2.4
r232 54 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=3.245
+ $X2=13.14 $Y2=3.33
r233 54 59 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=13.14 $Y=3.245
+ $X2=13.14 $Y2=2.4
r234 50 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.045 $Y=3.245
+ $X2=12.045 $Y2=3.33
r235 50 52 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=12.045 $Y=3.245
+ $X2=12.045 $Y2=2.805
r236 46 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.46 $Y=3.245
+ $X2=8.46 $Y2=3.33
r237 46 48 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=8.46 $Y=3.245
+ $X2=8.46 $Y2=2.475
r238 42 132 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.42 $Y=3.245
+ $X2=7.42 $Y2=3.33
r239 42 44 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=7.42 $Y=3.245
+ $X2=7.42 $Y2=2.795
r240 38 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=3.245
+ $X2=5.16 $Y2=3.33
r241 38 40 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.16 $Y=3.245
+ $X2=5.16 $Y2=2.81
r242 37 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.075 $Y2=3.33
r243 36 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=3.33
+ $X2=5.16 $Y2=3.33
r244 36 37 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.995 $Y=3.33
+ $X2=4.24 $Y2=3.33
r245 32 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=3.245
+ $X2=4.075 $Y2=3.33
r246 32 34 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.075 $Y=3.245
+ $X2=4.075 $Y2=2.81
r247 28 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r248 28 30 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.805
r249 9 59 300 $w=1.7e-07 $l=3.79737e-07 $layer=licon1_PDIFF $count=2 $X=12.905
+ $Y=2.12 $X2=13.14 $Y2=2.4
r250 9 56 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=12.905
+ $Y=2.12 $X2=13.14 $Y2=1.985
r251 8 52 600 $w=1.7e-07 $l=3.51034e-07 $layer=licon1_PDIFF $count=1 $X=11.845
+ $Y=2.54 $X2=12.045 $Y2=2.805
r252 7 138 600 $w=1.7e-07 $l=3.995e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=2.54 $X2=10.905 $Y2=2.815
r253 6 48 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.325
+ $Y=1.96 $X2=8.46 $Y2=2.475
r254 5 44 600 $w=1.7e-07 $l=3.21364e-07 $layer=licon1_PDIFF $count=1 $X=7.31
+ $Y=2.54 $X2=7.46 $Y2=2.795
r255 4 40 600 $w=1.7e-07 $l=1.03998e-06 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=1.84 $X2=5.16 $Y2=2.81
r256 3 34 600 $w=1.7e-07 $l=1.03998e-06 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=1.84 $X2=4.075 $Y2=2.81
r257 2 61 600 $w=1.7e-07 $l=8.44364e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=2.32 $X2=2.98 $Y2=3.055
r258 1 30 600 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.32 $X2=0.73 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%A_284_464# 1 2 3 4 5 18 22 25 26 27 28 29
+ 30 33 35 36 37 38 42 46 49 50 55 56
c156 56 0 1.90908e-19 $X=3.99 $Y=2.387
c157 38 0 1.32863e-19 $X=6.005 $Y=2.39
r158 49 50 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=2.795
+ $X2=2.22 $Y2=2.795
r159 44 46 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=6.13 $Y=2.475
+ $X2=6.13 $Y2=2.75
r160 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.03 $Y=0.7
+ $X2=6.03 $Y2=0.865
r161 39 56 5.10356 $w=1.72e-07 $l=8.6487e-08 $layer=LI1_cond $X=4.075 $Y=2.39
+ $X2=3.99 $Y2=2.387
r162 38 44 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.005 $Y=2.39
+ $X2=6.13 $Y2=2.475
r163 38 39 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=6.005 $Y=2.39
+ $X2=4.075 $Y2=2.39
r164 36 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.905 $Y=0.615
+ $X2=6.03 $Y2=0.7
r165 36 37 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=5.905 $Y=0.615
+ $X2=4.075 $Y2=0.615
r166 35 56 1.39518 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=3.99 $Y=2.3 $X2=3.99
+ $Y2=2.387
r167 34 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.185
+ $X2=3.99 $Y2=1.1
r168 34 35 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=3.99 $Y=1.185
+ $X2=3.99 $Y2=2.3
r169 33 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.015
+ $X2=3.99 $Y2=1.1
r170 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.99 $Y=0.7
+ $X2=4.075 $Y2=0.615
r171 32 33 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.99 $Y=0.7
+ $X2=3.99 $Y2=1.015
r172 31 52 4.16448 $w=1.75e-07 $l=1.25e-07 $layer=LI1_cond $X=3.68 $Y=2.387
+ $X2=3.555 $Y2=2.387
r173 30 56 5.10356 $w=1.72e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=2.387
+ $X2=3.99 $Y2=2.387
r174 30 31 14.2597 $w=1.73e-07 $l=2.25e-07 $layer=LI1_cond $X=3.905 $Y=2.387
+ $X2=3.68 $Y2=2.387
r175 29 54 3.20527 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=3.555 $Y=2.63
+ $X2=3.555 $Y2=2.805
r176 28 52 2.93179 $w=2.5e-07 $l=8.8e-08 $layer=LI1_cond $X=3.555 $Y=2.475
+ $X2=3.555 $Y2=2.387
r177 28 29 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=3.555 $Y=2.475
+ $X2=3.555 $Y2=2.63
r178 26 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=1.1
+ $X2=3.99 $Y2=1.1
r179 26 27 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=3.905 $Y=1.1
+ $X2=2.89 $Y2=1.1
r180 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.805 $Y=1.015
+ $X2=2.89 $Y2=1.1
r181 24 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.805 $Y=0.765
+ $X2=2.805 $Y2=1.015
r182 22 54 3.9379 $w=1.7e-07 $l=1.63936e-07 $layer=LI1_cond $X=3.43 $Y=2.715
+ $X2=3.555 $Y2=2.805
r183 22 50 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.43 $Y=2.715
+ $X2=2.22 $Y2=2.715
r184 18 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=0.68
+ $X2=2.805 $Y2=0.765
r185 18 20 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.72 $Y=0.68
+ $X2=2.26 $Y2=0.68
r186 5 46 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=6.025
+ $Y=2.54 $X2=6.17 $Y2=2.75
r187 4 54 600 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=2.32 $X2=3.515 $Y2=2.815
r188 4 52 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=2.32 $X2=3.515 $Y2=2.465
r189 3 49 300 $w=1.7e-07 $l=8.39553e-07 $layer=licon1_PDIFF $count=2 $X=1.42
+ $Y=2.32 $X2=2.055 $Y2=2.795
r190 2 42 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.925
+ $Y=0.655 $X2=6.07 $Y2=0.865
r191 1 20 182 $w=1.7e-07 $l=3.94208e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.405 $X2=2.26 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%Q 1 2 7 8 9 10 11 12 13
r13 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=2.405
+ $X2=13.64 $Y2=2.775
r14 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=13.64 $Y=1.985
+ $X2=13.64 $Y2=2.405
r15 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=13.64 $Y=1.665
+ $X2=13.64 $Y2=1.985
r16 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=1.295
+ $X2=13.64 $Y2=1.665
r17 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=0.925
+ $X2=13.64 $Y2=1.295
r18 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.64 $Y=0.515
+ $X2=13.64 $Y2=0.925
r19 2 13 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=13.485
+ $Y=1.84 $X2=13.64 $Y2=2.815
r20 2 11 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=13.485
+ $Y=1.84 $X2=13.64 $Y2=1.985
r21 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.5
+ $Y=0.37 $X2=13.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%VGND 1 2 3 4 5 6 21 25 29 33 37 39 49 54 59
+ 64 74 75 78 83 86 89 95 98 101
r118 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r119 98 99 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r120 95 96 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r121 89 92 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=4.985 $Y=0
+ $X2=4.985 $Y2=0.275
r122 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r123 85 86 10.9331 $w=4.43e-07 $l=2.45e-07 $layer=LI1_cond $X=3.82 $Y=0.137
+ $X2=4.065 $Y2=0.137
r124 81 85 5.69747 $w=4.43e-07 $l=2.2e-07 $layer=LI1_cond $X=3.6 $Y=0.137
+ $X2=3.82 $Y2=0.137
r125 81 83 5.23558 $w=4.43e-07 $l=2.5e-08 $layer=LI1_cond $X=3.6 $Y=0.137
+ $X2=3.575 $Y2=0.137
r126 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r127 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r128 75 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r129 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r130 72 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.14 $Y2=0
r131 72 74 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.68 $Y2=0
r132 71 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r133 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r134 68 71 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r135 68 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r136 67 70 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r137 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r138 65 98 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=11.2 $Y=0 $X2=10.965
+ $Y2=0
r139 65 67 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=11.2 $Y=0 $X2=11.28
+ $Y2=0
r140 64 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=13.14 $Y2=0
r141 64 70 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=12.72 $Y2=0
r142 63 99 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r143 63 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r144 62 63 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r145 60 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.22 $Y=0 $X2=8.055
+ $Y2=0
r146 60 62 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.22 $Y=0 $X2=8.4
+ $Y2=0
r147 59 98 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=10.73 $Y=0
+ $X2=10.965 $Y2=0
r148 59 62 152.011 $w=1.68e-07 $l=2.33e-06 $layer=LI1_cond $X=10.73 $Y=0 $X2=8.4
+ $Y2=0
r149 58 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r150 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r151 55 89 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=4.985
+ $Y2=0
r152 55 57 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r153 54 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.89 $Y=0 $X2=8.055
+ $Y2=0
r154 54 57 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=7.89 $Y=0 $X2=5.52
+ $Y2=0
r155 53 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r156 53 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r157 52 86 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.56 $Y=0
+ $X2=4.065 $Y2=0
r158 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r159 49 89 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.985
+ $Y2=0
r160 49 52 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.56
+ $Y2=0
r161 48 82 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r162 48 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r163 47 83 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=1.2 $Y=0
+ $X2=3.575 $Y2=0
r164 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r165 45 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r166 45 47 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r167 42 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r168 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r169 39 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r170 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r171 37 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r172 37 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.52 $Y2=0
r173 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.14 $Y=0.555
+ $X2=13.14 $Y2=0.965
r174 31 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0
r175 31 33 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0.555
r176 27 98 1.91284 $w=4.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.965 $Y=0.085
+ $X2=10.965 $Y2=0
r177 27 29 10.9428 $w=4.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.965 $Y=0.085
+ $X2=10.965 $Y2=0.515
r178 23 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.055 $Y=0.085
+ $X2=8.055 $Y2=0
r179 23 25 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.055 $Y=0.085
+ $X2=8.055 $Y2=0.535
r180 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r181 19 21 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.65
r182 6 35 182 $w=1.7e-07 $l=7.25655e-07 $layer=licon1_NDIFF $count=1 $X=12.92
+ $Y=0.37 $X2=13.21 $Y2=0.965
r183 6 33 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=12.92
+ $Y=0.37 $X2=13.14 $Y2=0.555
r184 5 29 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=10.765
+ $Y=0.37 $X2=10.965 $Y2=0.515
r185 4 25 182 $w=1.7e-07 $l=2.73496e-07 $layer=licon1_NDIFF $count=1 $X=7.835
+ $Y=0.655 $X2=8.055 $Y2=0.535
r186 3 92 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.135 $X2=4.985 $Y2=0.275
r187 2 85 182 $w=1.7e-07 $l=3.59166e-07 $layer=licon1_NDIFF $count=1 $X=3.52
+ $Y=0.405 $X2=3.82 $Y2=0.275
r188 1 21 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.44 $X2=0.78 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTN_1%noxref_24 1 2 9 11 12 15
r37 13 15 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.225 $Y=0.425
+ $X2=3.225 $Y2=0.615
r38 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=3.225 $Y2=0.425
r39 11 12 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=1.495 $Y2=0.34
r40 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.33 $Y=0.425
+ $X2=1.495 $Y2=0.34
r41 7 9 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.33 $Y=0.425 $X2=1.33
+ $Y2=0.575
r42 2 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.08
+ $Y=0.405 $X2=3.225 $Y2=0.615
r43 1 9 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.405 $X2=1.33 $Y2=0.575
.ends

