* File: sky130_fd_sc_hs__ebufn_4.pxi.spice
* Created: Thu Aug 27 20:44:10 2020
* 
x_PM_SKY130_FD_SC_HS__EBUFN_4%A N_A_c_124_n N_A_M1012_g N_A_M1003_g A
+ PM_SKY130_FD_SC_HS__EBUFN_4%A
x_PM_SKY130_FD_SC_HS__EBUFN_4%A_208_74# N_A_208_74#_M1011_d N_A_208_74#_M1015_d
+ N_A_208_74#_c_158_n N_A_208_74#_c_159_n N_A_208_74#_c_160_n
+ N_A_208_74#_M1006_g N_A_208_74#_c_161_n N_A_208_74#_c_162_n
+ N_A_208_74#_M1007_g N_A_208_74#_c_163_n N_A_208_74#_c_164_n
+ N_A_208_74#_M1009_g N_A_208_74#_c_165_n N_A_208_74#_c_166_n
+ N_A_208_74#_M1017_g N_A_208_74#_c_167_n N_A_208_74#_c_168_n
+ N_A_208_74#_c_169_n N_A_208_74#_c_174_n N_A_208_74#_c_173_n
+ N_A_208_74#_c_170_n N_A_208_74#_c_171_n N_A_208_74#_c_172_n
+ PM_SKY130_FD_SC_HS__EBUFN_4%A_208_74#
x_PM_SKY130_FD_SC_HS__EBUFN_4%TE_B N_TE_B_M1011_g N_TE_B_c_267_n N_TE_B_c_279_n
+ N_TE_B_M1015_g N_TE_B_c_268_n N_TE_B_c_281_n N_TE_B_M1000_g N_TE_B_c_269_n
+ N_TE_B_c_283_n N_TE_B_M1001_g N_TE_B_c_270_n N_TE_B_c_285_n N_TE_B_M1002_g
+ N_TE_B_c_271_n N_TE_B_c_287_n N_TE_B_M1018_g N_TE_B_c_272_n N_TE_B_c_273_n
+ N_TE_B_c_274_n N_TE_B_c_275_n TE_B N_TE_B_c_277_n N_TE_B_c_278_n
+ PM_SKY130_FD_SC_HS__EBUFN_4%TE_B
x_PM_SKY130_FD_SC_HS__EBUFN_4%A_27_368# N_A_27_368#_M1003_s N_A_27_368#_M1012_s
+ N_A_27_368#_c_410_n N_A_27_368#_M1004_g N_A_27_368#_M1005_g
+ N_A_27_368#_c_411_n N_A_27_368#_M1008_g N_A_27_368#_M1013_g
+ N_A_27_368#_c_412_n N_A_27_368#_M1010_g N_A_27_368#_M1014_g
+ N_A_27_368#_c_413_n N_A_27_368#_M1016_g N_A_27_368#_M1019_g
+ N_A_27_368#_c_403_n N_A_27_368#_c_414_n N_A_27_368#_c_415_n
+ N_A_27_368#_c_416_n N_A_27_368#_c_417_n N_A_27_368#_c_418_n
+ N_A_27_368#_c_419_n N_A_27_368#_c_420_n N_A_27_368#_c_421_n
+ N_A_27_368#_c_404_n N_A_27_368#_c_405_n N_A_27_368#_c_518_p
+ N_A_27_368#_c_406_n N_A_27_368#_c_407_n N_A_27_368#_c_423_n
+ N_A_27_368#_c_408_n N_A_27_368#_c_409_n PM_SKY130_FD_SC_HS__EBUFN_4%A_27_368#
x_PM_SKY130_FD_SC_HS__EBUFN_4%VPWR N_VPWR_M1012_d N_VPWR_M1000_s N_VPWR_M1002_s
+ N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_572_n N_VPWR_c_573_n
+ N_VPWR_c_574_n VPWR N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_568_n
+ N_VPWR_c_578_n N_VPWR_c_579_n PM_SKY130_FD_SC_HS__EBUFN_4%VPWR
x_PM_SKY130_FD_SC_HS__EBUFN_4%A_348_368# N_A_348_368#_M1000_d
+ N_A_348_368#_M1001_d N_A_348_368#_M1018_d N_A_348_368#_M1008_s
+ N_A_348_368#_M1016_s N_A_348_368#_c_652_n N_A_348_368#_c_642_n
+ N_A_348_368#_c_658_n N_A_348_368#_c_643_n N_A_348_368#_c_644_n
+ N_A_348_368#_c_645_n N_A_348_368#_c_669_n N_A_348_368#_c_646_n
+ N_A_348_368#_c_647_n N_A_348_368#_c_722_p N_A_348_368#_c_648_n
+ N_A_348_368#_c_649_n N_A_348_368#_c_672_n N_A_348_368#_c_713_n
+ N_A_348_368#_c_650_n PM_SKY130_FD_SC_HS__EBUFN_4%A_348_368#
x_PM_SKY130_FD_SC_HS__EBUFN_4%Z N_Z_M1005_s N_Z_M1014_s N_Z_M1004_d N_Z_M1010_d
+ N_Z_c_730_n N_Z_c_734_n N_Z_c_742_n N_Z_c_731_n N_Z_c_726_n N_Z_c_727_n
+ N_Z_c_757_n N_Z_c_728_n N_Z_c_729_n Z Z Z PM_SKY130_FD_SC_HS__EBUFN_4%Z
x_PM_SKY130_FD_SC_HS__EBUFN_4%VGND N_VGND_M1003_d N_VGND_M1006_d N_VGND_M1009_d
+ N_VGND_c_794_n N_VGND_c_795_n N_VGND_c_796_n N_VGND_c_797_n N_VGND_c_798_n
+ N_VGND_c_799_n N_VGND_c_800_n VGND N_VGND_c_801_n N_VGND_c_802_n
+ N_VGND_c_803_n N_VGND_c_804_n PM_SKY130_FD_SC_HS__EBUFN_4%VGND
x_PM_SKY130_FD_SC_HS__EBUFN_4%A_378_74# N_A_378_74#_M1006_s N_A_378_74#_M1007_s
+ N_A_378_74#_M1017_s N_A_378_74#_M1013_d N_A_378_74#_M1019_d
+ N_A_378_74#_c_866_n N_A_378_74#_c_867_n N_A_378_74#_c_868_n
+ N_A_378_74#_c_869_n N_A_378_74#_c_870_n N_A_378_74#_c_896_n
+ N_A_378_74#_c_871_n N_A_378_74#_c_872_n N_A_378_74#_c_923_n
+ N_A_378_74#_c_873_n N_A_378_74#_c_874_n N_A_378_74#_c_875_n
+ N_A_378_74#_c_876_n PM_SKY130_FD_SC_HS__EBUFN_4%A_378_74#
cc_1 VNB N_A_c_124_n 0.0358282f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_M1003_g 0.0263754f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.74
cc_3 VNB A 0.00396202f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_208_74#_c_158_n 0.0205453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_208_74#_c_159_n 0.011951f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_6 VNB N_A_208_74#_c_160_n 0.0166173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_208_74#_c_161_n 0.0122721f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_8 VNB N_A_208_74#_c_162_n 0.01433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_208_74#_c_163_n 0.0122636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_208_74#_c_164_n 0.0143385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_208_74#_c_165_n 0.0200371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_208_74#_c_166_n 0.0146143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_208_74#_c_167_n 0.00514785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_208_74#_c_168_n 0.00511446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_208_74#_c_169_n 0.00511446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_208_74#_c_170_n 0.00848374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_208_74#_c_171_n 0.00568136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_208_74#_c_172_n 0.0754207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_TE_B_c_267_n 0.014558f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.74
cc_20 VNB N_TE_B_c_268_n 0.0209237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_TE_B_c_269_n 0.00646238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_TE_B_c_270_n 0.00552156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_TE_B_c_271_n 0.0103914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_TE_B_c_272_n 0.00469483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_TE_B_c_273_n 0.00489103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_TE_B_c_274_n 0.0036966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_TE_B_c_275_n 0.0036966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB TE_B 0.00702428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_TE_B_c_277_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_TE_B_c_278_n 0.0192479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_368#_M1005_g 0.0214935f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_32 VNB N_A_27_368#_M1013_g 0.0209312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_368#_M1014_g 0.0211723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_368#_M1019_g 0.0285164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_368#_c_403_n 0.0280304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_368#_c_404_n 0.0025686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_368#_c_405_n 0.00606935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_368#_c_406_n 0.0112533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_368#_c_407_n 0.0248753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_368#_c_408_n 0.0135381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_368#_c_409_n 0.114625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_568_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Z_c_726_n 0.00225436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Z_c_727_n 0.00229628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Z_c_728_n 0.00122079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Z_c_729_n 0.00176823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_794_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_48 VNB N_VGND_c_795_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_796_n 0.00452091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_797_n 0.0363752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_798_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_799_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_800_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_801_n 0.018117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_802_n 0.0569796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_803_n 0.328933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_804_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_378_74#_c_866_n 0.00221841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_378_74#_c_867_n 0.0063992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_378_74#_c_868_n 2.51175e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_378_74#_c_869_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_378_74#_c_870_n 0.00578259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_378_74#_c_871_n 0.0027626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_378_74#_c_872_n 0.00163793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_378_74#_c_873_n 0.0122413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_378_74#_c_874_n 0.0364928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_378_74#_c_875_n 7.52762e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_378_74#_c_876_n 0.00121874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VPB N_A_c_124_n 0.0256832f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_70 VPB A 0.00486006f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_71 VPB N_A_208_74#_c_173_n 0.00533118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_TE_B_c_279_n 0.0198654f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.74
cc_73 VPB N_TE_B_c_268_n 0.026733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_TE_B_c_281_n 0.0191931f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.465
cc_75 VPB N_TE_B_c_269_n 0.00891526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_TE_B_c_283_n 0.01477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_TE_B_c_270_n 0.00810834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_TE_B_c_285_n 0.0148977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_TE_B_c_271_n 0.0129907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_TE_B_c_287_n 0.0151359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_TE_B_c_272_n 0.0122435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_TE_B_c_273_n 0.00437671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_TE_B_c_274_n 0.00410577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_TE_B_c_275_n 0.00402089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_27_368#_c_410_n 0.0148126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_27_368#_c_411_n 0.0144924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_27_368#_c_412_n 0.0144924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_27_368#_c_413_n 0.0180496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_368#_c_414_n 0.00536733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_27_368#_c_415_n 0.0114247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_27_368#_c_416_n 0.0187408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_368#_c_417_n 0.0091553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_368#_c_418_n 0.00469589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_27_368#_c_419_n 0.00513674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_27_368#_c_420_n 0.0034565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_368#_c_421_n 0.00108034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_368#_c_407_n 0.0127952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_27_368#_c_423_n 0.00723806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_27_368#_c_409_n 0.0292369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_569_n 0.00396699f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.465
cc_101 VPB N_VPWR_c_570_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_571_n 0.0157448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_572_n 0.00471226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_573_n 0.0377381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_574_n 0.00601619f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_575_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_576_n 0.0591189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_568_n 0.0823537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_578_n 0.00647446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_579_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_348_368#_c_642_n 0.00114639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_348_368#_c_643_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_348_368#_c_644_n 0.00212406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_348_368#_c_645_n 0.00217419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_348_368#_c_646_n 0.0028338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_348_368#_c_647_n 0.00171072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_348_368#_c_648_n 0.0122025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_348_368#_c_649_n 0.0503972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_348_368#_c_650_n 0.00167433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_Z_c_730_n 0.00183525f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.54
cc_121 VPB N_Z_c_731_n 0.00179576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_Z_c_728_n 0.0010334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB Z 0.00133625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 N_A_c_124_n N_A_208_74#_c_174_n 0.00111598f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_c_124_n N_A_208_74#_c_173_n 5.55952e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_126 A N_A_208_74#_c_173_n 0.003836f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_127 A N_A_208_74#_c_170_n 0.0049962f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A_c_124_n N_TE_B_c_279_n 0.0364083f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_c_124_n N_TE_B_c_272_n 0.00548243f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_c_124_n TE_B 2.12581e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_M1003_g TE_B 6.22691e-19 $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_132 A TE_B 0.0199149f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A_c_124_n N_TE_B_c_277_n 0.0206413f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_134 A N_TE_B_c_277_n 0.00464778f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A_M1003_g N_TE_B_c_278_n 0.0159419f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_M1003_g N_A_27_368#_c_403_n 0.00241184f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_c_124_n N_A_27_368#_c_414_n 5.30183e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_c_124_n N_A_27_368#_c_416_n 0.00494922f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A_c_124_n N_A_27_368#_c_417_n 0.0117611f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_140 A N_A_27_368#_c_417_n 0.0103329f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_141 N_A_c_124_n N_A_27_368#_c_406_n 0.00239983f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_c_124_n N_A_27_368#_c_407_n 0.0150151f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_M1003_g N_A_27_368#_c_407_n 0.0039401f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_144 A N_A_27_368#_c_407_n 0.0365496f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_145 N_A_c_124_n N_VPWR_c_569_n 0.00947766f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_c_124_n N_VPWR_c_575_n 0.00413917f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_c_124_n N_VPWR_c_568_n 0.00402136f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_c_124_n N_VGND_c_794_n 0.00129795f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_M1003_g N_VGND_c_794_n 0.0144322f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_150 A N_VGND_c_794_n 0.01106f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A_M1003_g N_VGND_c_801_n 0.00383152f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_M1003_g N_VGND_c_803_n 0.00761327f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_208_74#_c_170_n N_TE_B_c_267_n 6.8085e-19 $X=1.615 $Y=1.145 $X2=0
+ $Y2=0
cc_154 N_A_208_74#_c_174_n N_TE_B_c_279_n 0.00658052f $X=1.205 $Y=2.02 $X2=0
+ $Y2=0
cc_155 N_A_208_74#_c_173_n N_TE_B_c_279_n 0.00412409f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_156 N_A_208_74#_c_159_n N_TE_B_c_268_n 0.0167668f $X=1.78 $Y=1.26 $X2=0 $Y2=0
cc_157 N_A_208_74#_c_173_n N_TE_B_c_268_n 0.0173987f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_158 N_A_208_74#_c_170_n N_TE_B_c_268_n 0.0163685f $X=1.615 $Y=1.145 $X2=0
+ $Y2=0
cc_159 N_A_208_74#_c_171_n N_TE_B_c_268_n 0.0046517f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_160 N_A_208_74#_c_173_n N_TE_B_c_281_n 0.00283047f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_161 N_A_208_74#_c_167_n N_TE_B_c_269_n 0.0167668f $X=2.245 $Y=1.26 $X2=0
+ $Y2=0
cc_162 N_A_208_74#_c_168_n N_TE_B_c_270_n 0.0167668f $X=2.675 $Y=1.26 $X2=0
+ $Y2=0
cc_163 N_A_208_74#_c_169_n N_TE_B_c_271_n 0.0167668f $X=3.105 $Y=1.26 $X2=0
+ $Y2=0
cc_164 N_A_208_74#_c_174_n N_TE_B_c_272_n 0.00108213f $X=1.205 $Y=2.02 $X2=0
+ $Y2=0
cc_165 N_A_208_74#_c_173_n N_TE_B_c_272_n 0.00757366f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_166 N_A_208_74#_c_158_n N_TE_B_c_273_n 0.0167668f $X=2.17 $Y=1.26 $X2=0 $Y2=0
cc_167 N_A_208_74#_c_173_n N_TE_B_c_273_n 9.62687e-19 $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_168 N_A_208_74#_c_161_n N_TE_B_c_274_n 0.0167668f $X=2.6 $Y=1.26 $X2=0 $Y2=0
cc_169 N_A_208_74#_c_163_n N_TE_B_c_275_n 0.0167668f $X=3.03 $Y=1.26 $X2=0 $Y2=0
cc_170 N_A_208_74#_c_173_n TE_B 0.0178111f $X=1.615 $Y=1.72 $X2=0 $Y2=0
cc_171 N_A_208_74#_c_170_n TE_B 0.0298967f $X=1.615 $Y=1.145 $X2=0 $Y2=0
cc_172 N_A_208_74#_c_171_n TE_B 0.0164997f $X=1.615 $Y=0.465 $X2=0 $Y2=0
cc_173 N_A_208_74#_c_172_n TE_B 0.00107199f $X=1.615 $Y=0.465 $X2=0 $Y2=0
cc_174 N_A_208_74#_c_159_n N_TE_B_c_277_n 0.00761709f $X=1.78 $Y=1.26 $X2=0
+ $Y2=0
cc_175 N_A_208_74#_c_170_n N_TE_B_c_277_n 0.00152275f $X=1.615 $Y=1.145 $X2=0
+ $Y2=0
cc_176 N_A_208_74#_c_171_n N_TE_B_c_277_n 0.00101764f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_177 N_A_208_74#_c_170_n N_TE_B_c_278_n 9.11108e-19 $X=1.615 $Y=1.145 $X2=0
+ $Y2=0
cc_178 N_A_208_74#_c_171_n N_TE_B_c_278_n 6.76457e-19 $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_179 N_A_208_74#_c_172_n N_TE_B_c_278_n 0.016396f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_180 N_A_208_74#_c_166_n N_A_27_368#_M1005_g 0.0193926f $X=3.535 $Y=1.185
+ $X2=0 $Y2=0
cc_181 N_A_208_74#_c_174_n N_A_27_368#_c_414_n 0.00673641f $X=1.205 $Y=2.02
+ $X2=0 $Y2=0
cc_182 N_A_208_74#_M1015_d N_A_27_368#_c_417_n 0.00829457f $X=1.055 $Y=1.84
+ $X2=0 $Y2=0
cc_183 N_A_208_74#_c_174_n N_A_27_368#_c_417_n 0.0145977f $X=1.205 $Y=2.02 $X2=0
+ $Y2=0
cc_184 N_A_208_74#_c_173_n N_A_27_368#_c_417_n 0.00592951f $X=1.615 $Y=1.72
+ $X2=0 $Y2=0
cc_185 N_A_208_74#_c_173_n N_A_27_368#_c_419_n 0.0107872f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_186 N_A_208_74#_c_174_n N_A_27_368#_c_420_n 0.0136474f $X=1.205 $Y=2.02 $X2=0
+ $Y2=0
cc_187 N_A_208_74#_c_173_n N_A_27_368#_c_420_n 0.0139991f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_188 N_A_208_74#_c_173_n N_A_27_368#_c_421_n 0.0057474f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_189 N_A_208_74#_c_170_n N_A_27_368#_c_421_n 0.00178624f $X=1.615 $Y=1.145
+ $X2=0 $Y2=0
cc_190 N_A_208_74#_c_161_n N_A_27_368#_c_404_n 0.00115704f $X=2.6 $Y=1.26 $X2=0
+ $Y2=0
cc_191 N_A_208_74#_c_170_n N_A_27_368#_c_404_n 0.00569129f $X=1.615 $Y=1.145
+ $X2=0 $Y2=0
cc_192 N_A_208_74#_c_161_n N_A_27_368#_c_408_n 0.00936976f $X=2.6 $Y=1.26 $X2=0
+ $Y2=0
cc_193 N_A_208_74#_c_165_n N_A_27_368#_c_409_n 0.0010213f $X=3.46 $Y=1.26 $X2=0
+ $Y2=0
cc_194 N_A_208_74#_c_173_n N_A_348_368#_M1000_d 0.00112287f $X=1.615 $Y=1.72
+ $X2=-0.19 $Y2=-0.245
cc_195 N_A_208_74#_c_171_n N_VGND_c_794_n 0.0285331f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_196 N_A_208_74#_c_172_n N_VGND_c_794_n 4.72719e-19 $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_197 N_A_208_74#_c_160_n N_VGND_c_795_n 0.0122493f $X=2.245 $Y=1.185 $X2=0
+ $Y2=0
cc_198 N_A_208_74#_c_161_n N_VGND_c_795_n 7.11061e-19 $X=2.6 $Y=1.26 $X2=0 $Y2=0
cc_199 N_A_208_74#_c_162_n N_VGND_c_795_n 0.0106722f $X=2.675 $Y=1.185 $X2=0
+ $Y2=0
cc_200 N_A_208_74#_c_164_n N_VGND_c_795_n 5.10431e-19 $X=3.105 $Y=1.185 $X2=0
+ $Y2=0
cc_201 N_A_208_74#_c_171_n N_VGND_c_795_n 0.00156286f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_202 N_A_208_74#_c_172_n N_VGND_c_795_n 3.15165e-19 $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_203 N_A_208_74#_c_162_n N_VGND_c_796_n 4.64001e-19 $X=2.675 $Y=1.185 $X2=0
+ $Y2=0
cc_204 N_A_208_74#_c_164_n N_VGND_c_796_n 0.0093975f $X=3.105 $Y=1.185 $X2=0
+ $Y2=0
cc_205 N_A_208_74#_c_166_n N_VGND_c_796_n 0.00154624f $X=3.535 $Y=1.185 $X2=0
+ $Y2=0
cc_206 N_A_208_74#_c_160_n N_VGND_c_797_n 0.00383152f $X=2.245 $Y=1.185 $X2=0
+ $Y2=0
cc_207 N_A_208_74#_c_171_n N_VGND_c_797_n 0.0367749f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_208 N_A_208_74#_c_172_n N_VGND_c_797_n 0.00827872f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_209 N_A_208_74#_c_162_n N_VGND_c_799_n 0.00383152f $X=2.675 $Y=1.185 $X2=0
+ $Y2=0
cc_210 N_A_208_74#_c_164_n N_VGND_c_799_n 0.00383152f $X=3.105 $Y=1.185 $X2=0
+ $Y2=0
cc_211 N_A_208_74#_c_166_n N_VGND_c_802_n 0.00430908f $X=3.535 $Y=1.185 $X2=0
+ $Y2=0
cc_212 N_A_208_74#_c_160_n N_VGND_c_803_n 0.00762539f $X=2.245 $Y=1.185 $X2=0
+ $Y2=0
cc_213 N_A_208_74#_c_162_n N_VGND_c_803_n 0.0075754f $X=2.675 $Y=1.185 $X2=0
+ $Y2=0
cc_214 N_A_208_74#_c_164_n N_VGND_c_803_n 0.0075754f $X=3.105 $Y=1.185 $X2=0
+ $Y2=0
cc_215 N_A_208_74#_c_166_n N_VGND_c_803_n 0.0081578f $X=3.535 $Y=1.185 $X2=0
+ $Y2=0
cc_216 N_A_208_74#_c_171_n N_VGND_c_803_n 0.0256312f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_217 N_A_208_74#_c_172_n N_VGND_c_803_n 0.0115893f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_218 N_A_208_74#_c_160_n N_A_378_74#_c_866_n 0.00122164f $X=2.245 $Y=1.185
+ $X2=0 $Y2=0
cc_219 N_A_208_74#_c_170_n N_A_378_74#_c_866_n 0.00957786f $X=1.615 $Y=1.145
+ $X2=0 $Y2=0
cc_220 N_A_208_74#_c_171_n N_A_378_74#_c_866_n 0.0518232f $X=1.615 $Y=0.465
+ $X2=0 $Y2=0
cc_221 N_A_208_74#_c_172_n N_A_378_74#_c_866_n 0.00601712f $X=1.615 $Y=0.465
+ $X2=0 $Y2=0
cc_222 N_A_208_74#_c_158_n N_A_378_74#_c_867_n 0.00129279f $X=2.17 $Y=1.26 $X2=0
+ $Y2=0
cc_223 N_A_208_74#_c_160_n N_A_378_74#_c_867_n 0.00749872f $X=2.245 $Y=1.185
+ $X2=0 $Y2=0
cc_224 N_A_208_74#_c_161_n N_A_378_74#_c_867_n 0.00643581f $X=2.6 $Y=1.26 $X2=0
+ $Y2=0
cc_225 N_A_208_74#_c_162_n N_A_378_74#_c_867_n 0.00721311f $X=2.675 $Y=1.185
+ $X2=0 $Y2=0
cc_226 N_A_208_74#_c_163_n N_A_378_74#_c_867_n 0.00129486f $X=3.03 $Y=1.26 $X2=0
+ $Y2=0
cc_227 N_A_208_74#_c_167_n N_A_378_74#_c_867_n 0.00365884f $X=2.245 $Y=1.26
+ $X2=0 $Y2=0
cc_228 N_A_208_74#_c_168_n N_A_378_74#_c_867_n 0.00251095f $X=2.675 $Y=1.26
+ $X2=0 $Y2=0
cc_229 N_A_208_74#_c_158_n N_A_378_74#_c_868_n 0.0096098f $X=2.17 $Y=1.26 $X2=0
+ $Y2=0
cc_230 N_A_208_74#_c_170_n N_A_378_74#_c_868_n 0.0137054f $X=1.615 $Y=1.145
+ $X2=0 $Y2=0
cc_231 N_A_208_74#_c_172_n N_A_378_74#_c_868_n 3.76302e-19 $X=1.615 $Y=0.465
+ $X2=0 $Y2=0
cc_232 N_A_208_74#_c_162_n N_A_378_74#_c_869_n 0.00111248f $X=2.675 $Y=1.185
+ $X2=0 $Y2=0
cc_233 N_A_208_74#_c_164_n N_A_378_74#_c_869_n 3.92313e-19 $X=3.105 $Y=1.185
+ $X2=0 $Y2=0
cc_234 N_A_208_74#_c_164_n N_A_378_74#_c_870_n 0.0122885f $X=3.105 $Y=1.185
+ $X2=0 $Y2=0
cc_235 N_A_208_74#_c_165_n N_A_378_74#_c_870_n 0.0024802f $X=3.46 $Y=1.26 $X2=0
+ $Y2=0
cc_236 N_A_208_74#_c_166_n N_A_378_74#_c_870_n 0.0121337f $X=3.535 $Y=1.185
+ $X2=0 $Y2=0
cc_237 N_A_208_74#_c_164_n N_A_378_74#_c_896_n 5.78934e-19 $X=3.105 $Y=1.185
+ $X2=0 $Y2=0
cc_238 N_A_208_74#_c_166_n N_A_378_74#_c_896_n 0.00767715f $X=3.535 $Y=1.185
+ $X2=0 $Y2=0
cc_239 N_A_208_74#_c_166_n N_A_378_74#_c_872_n 0.00322875f $X=3.535 $Y=1.185
+ $X2=0 $Y2=0
cc_240 N_A_208_74#_c_163_n N_A_378_74#_c_875_n 0.0109545f $X=3.03 $Y=1.26 $X2=0
+ $Y2=0
cc_241 N_A_208_74#_c_164_n N_A_378_74#_c_875_n 9.32193e-19 $X=3.105 $Y=1.185
+ $X2=0 $Y2=0
cc_242 N_TE_B_c_287_n N_A_27_368#_c_410_n 0.010534f $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_243 N_TE_B_c_279_n N_A_27_368#_c_417_n 0.0177405f $X=0.98 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_TE_B_c_268_n N_A_27_368#_c_417_n 8.76722e-19 $X=2.02 $Y=1.65 $X2=0
+ $Y2=0
cc_245 N_TE_B_c_279_n N_A_27_368#_c_418_n 0.00424479f $X=0.98 $Y=1.765 $X2=0
+ $Y2=0
cc_246 N_TE_B_c_281_n N_A_27_368#_c_418_n 0.00398125f $X=2.11 $Y=1.765 $X2=0
+ $Y2=0
cc_247 N_TE_B_c_268_n N_A_27_368#_c_419_n 0.00710522f $X=2.02 $Y=1.65 $X2=0
+ $Y2=0
cc_248 N_TE_B_c_281_n N_A_27_368#_c_419_n 0.0166834f $X=2.11 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_TE_B_c_269_n N_A_27_368#_c_419_n 0.00395544f $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_250 N_TE_B_c_283_n N_A_27_368#_c_419_n 0.00476803f $X=2.56 $Y=1.765 $X2=0
+ $Y2=0
cc_251 N_TE_B_c_279_n N_A_27_368#_c_420_n 6.4739e-19 $X=0.98 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_TE_B_c_268_n N_A_27_368#_c_420_n 8.92373e-19 $X=2.02 $Y=1.65 $X2=0
+ $Y2=0
cc_253 N_TE_B_c_281_n N_A_27_368#_c_421_n 0.00475251f $X=2.11 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_TE_B_c_269_n N_A_27_368#_c_421_n 0.00504799f $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_255 N_TE_B_c_283_n N_A_27_368#_c_421_n 0.00588941f $X=2.56 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_TE_B_c_285_n N_A_27_368#_c_421_n 3.33195e-19 $X=3.01 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_TE_B_c_273_n N_A_27_368#_c_421_n 3.98382e-19 $X=2.11 $Y=1.67 $X2=0
+ $Y2=0
cc_258 N_TE_B_c_274_n N_A_27_368#_c_421_n 0.00507112f $X=2.56 $Y=1.67 $X2=0
+ $Y2=0
cc_259 N_TE_B_c_275_n N_A_27_368#_c_421_n 2.0327e-19 $X=3.01 $Y=1.67 $X2=0 $Y2=0
cc_260 N_TE_B_c_269_n N_A_27_368#_c_404_n 0.00346529f $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_261 N_TE_B_c_274_n N_A_27_368#_c_404_n 7.22911e-19 $X=2.56 $Y=1.67 $X2=0
+ $Y2=0
cc_262 N_TE_B_c_270_n N_A_27_368#_c_408_n 0.00658386f $X=2.92 $Y=1.65 $X2=0
+ $Y2=0
cc_263 N_TE_B_c_271_n N_A_27_368#_c_408_n 0.0104102f $X=3.37 $Y=1.65 $X2=0 $Y2=0
cc_264 N_TE_B_c_274_n N_A_27_368#_c_408_n 0.00658868f $X=2.56 $Y=1.67 $X2=0
+ $Y2=0
cc_265 N_TE_B_c_275_n N_A_27_368#_c_408_n 0.00444171f $X=3.01 $Y=1.67 $X2=0
+ $Y2=0
cc_266 N_TE_B_c_271_n N_A_27_368#_c_409_n 0.0102891f $X=3.37 $Y=1.65 $X2=0 $Y2=0
cc_267 N_TE_B_c_279_n N_VPWR_c_569_n 0.0175124f $X=0.98 $Y=1.765 $X2=0 $Y2=0
cc_268 N_TE_B_c_281_n N_VPWR_c_570_n 0.0143533f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_269 N_TE_B_c_283_n N_VPWR_c_570_n 0.00646001f $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_270 N_TE_B_c_285_n N_VPWR_c_570_n 3.99197e-19 $X=3.01 $Y=1.765 $X2=0 $Y2=0
cc_271 N_TE_B_c_283_n N_VPWR_c_571_n 0.00304555f $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_272 N_TE_B_c_285_n N_VPWR_c_571_n 0.00413917f $X=3.01 $Y=1.765 $X2=0 $Y2=0
cc_273 N_TE_B_c_283_n N_VPWR_c_572_n 4.52399e-19 $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_274 N_TE_B_c_285_n N_VPWR_c_572_n 0.0129243f $X=3.01 $Y=1.765 $X2=0 $Y2=0
cc_275 N_TE_B_c_287_n N_VPWR_c_572_n 0.00445463f $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_276 N_TE_B_c_279_n N_VPWR_c_573_n 0.00413917f $X=0.98 $Y=1.765 $X2=0 $Y2=0
cc_277 N_TE_B_c_281_n N_VPWR_c_573_n 0.00304555f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_278 N_TE_B_c_287_n N_VPWR_c_576_n 0.0044313f $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_279 N_TE_B_c_279_n N_VPWR_c_568_n 0.00403443f $X=0.98 $Y=1.765 $X2=0 $Y2=0
cc_280 N_TE_B_c_281_n N_VPWR_c_568_n 0.00401174f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_281 N_TE_B_c_283_n N_VPWR_c_568_n 0.00396372f $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_282 N_TE_B_c_285_n N_VPWR_c_568_n 0.00817726f $X=3.01 $Y=1.765 $X2=0 $Y2=0
cc_283 N_TE_B_c_287_n N_VPWR_c_568_n 0.00853445f $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_284 N_TE_B_c_281_n N_A_348_368#_c_652_n 0.0100509f $X=2.11 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_TE_B_c_269_n N_A_348_368#_c_652_n 3.64605e-19 $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_286 N_TE_B_c_283_n N_A_348_368#_c_652_n 0.0132117f $X=2.56 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_TE_B_c_270_n N_A_348_368#_c_652_n 5.64341e-19 $X=2.92 $Y=1.65 $X2=0
+ $Y2=0
cc_288 N_TE_B_c_283_n N_A_348_368#_c_642_n 7.30235e-19 $X=2.56 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_TE_B_c_270_n N_A_348_368#_c_642_n 0.00372332f $X=2.92 $Y=1.65 $X2=0
+ $Y2=0
cc_290 N_TE_B_c_283_n N_A_348_368#_c_658_n 0.00404286f $X=2.56 $Y=1.765 $X2=0
+ $Y2=0
cc_291 N_TE_B_c_285_n N_A_348_368#_c_658_n 0.00229356f $X=3.01 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_TE_B_c_283_n N_A_348_368#_c_643_n 0.00423981f $X=2.56 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_TE_B_c_285_n N_A_348_368#_c_643_n 0.00148725f $X=3.01 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_TE_B_c_270_n N_A_348_368#_c_644_n 0.0010235f $X=2.92 $Y=1.65 $X2=0
+ $Y2=0
cc_295 N_TE_B_c_285_n N_A_348_368#_c_644_n 0.0127103f $X=3.01 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_TE_B_c_271_n N_A_348_368#_c_644_n 0.00594793f $X=3.37 $Y=1.65 $X2=0
+ $Y2=0
cc_297 N_TE_B_c_287_n N_A_348_368#_c_644_n 0.0118656f $X=3.46 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_TE_B_c_275_n N_A_348_368#_c_644_n 6.89848e-19 $X=3.01 $Y=1.67 $X2=0
+ $Y2=0
cc_299 N_TE_B_c_271_n N_A_348_368#_c_645_n 3.61478e-19 $X=3.37 $Y=1.65 $X2=0
+ $Y2=0
cc_300 N_TE_B_c_287_n N_A_348_368#_c_645_n 6.17533e-19 $X=3.46 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_TE_B_c_285_n N_A_348_368#_c_669_n 7.24077e-19 $X=3.01 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_TE_B_c_287_n N_A_348_368#_c_669_n 0.0112031f $X=3.46 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_TE_B_c_287_n N_A_348_368#_c_647_n 0.0032261f $X=3.46 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_TE_B_c_281_n N_A_348_368#_c_672_n 0.00471362f $X=2.11 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_TE_B_c_287_n N_Z_c_734_n 2.48499e-19 $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_306 N_TE_B_c_278_n N_VGND_c_794_n 0.0133028f $X=1.065 $Y=1.22 $X2=0 $Y2=0
cc_307 N_TE_B_c_278_n N_VGND_c_797_n 0.00383152f $X=1.065 $Y=1.22 $X2=0 $Y2=0
cc_308 N_TE_B_c_278_n N_VGND_c_803_n 0.00762539f $X=1.065 $Y=1.22 $X2=0 $Y2=0
cc_309 N_TE_B_c_269_n N_A_378_74#_c_867_n 4.57305e-19 $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_310 N_TE_B_c_273_n N_A_378_74#_c_867_n 0.00157449f $X=2.11 $Y=1.67 $X2=0
+ $Y2=0
cc_311 N_TE_B_c_268_n N_A_378_74#_c_868_n 0.00111257f $X=2.02 $Y=1.65 $X2=0
+ $Y2=0
cc_312 N_TE_B_c_271_n N_A_378_74#_c_870_n 6.30494e-19 $X=3.37 $Y=1.65 $X2=0
+ $Y2=0
cc_313 N_TE_B_c_275_n N_A_378_74#_c_870_n 2.8721e-19 $X=3.01 $Y=1.67 $X2=0 $Y2=0
cc_314 N_A_27_368#_c_417_n N_VPWR_M1012_d 0.00721344f $X=1.46 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A_27_368#_c_419_n N_VPWR_M1000_s 0.00354253f $X=2.36 $Y=2.145 $X2=0
+ $Y2=0
cc_316 N_A_27_368#_c_421_n N_VPWR_M1000_s 0.00266592f $X=2.445 $Y=2.06 $X2=0
+ $Y2=0
cc_317 N_A_27_368#_c_416_n N_VPWR_c_569_n 0.0170312f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_318 N_A_27_368#_c_417_n N_VPWR_c_569_n 0.0186768f $X=1.46 $Y=2.475 $X2=0
+ $Y2=0
cc_319 N_A_27_368#_c_416_n N_VPWR_c_575_n 0.0124046f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_320 N_A_27_368#_c_410_n N_VPWR_c_576_n 0.00278271f $X=3.91 $Y=1.765 $X2=0
+ $Y2=0
cc_321 N_A_27_368#_c_411_n N_VPWR_c_576_n 0.00278271f $X=4.36 $Y=1.765 $X2=0
+ $Y2=0
cc_322 N_A_27_368#_c_412_n N_VPWR_c_576_n 0.00278271f $X=4.81 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A_27_368#_c_413_n N_VPWR_c_576_n 0.00278271f $X=5.26 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_A_27_368#_c_410_n N_VPWR_c_568_n 0.00353907f $X=3.91 $Y=1.765 $X2=0
+ $Y2=0
cc_325 N_A_27_368#_c_411_n N_VPWR_c_568_n 0.00353823f $X=4.36 $Y=1.765 $X2=0
+ $Y2=0
cc_326 N_A_27_368#_c_412_n N_VPWR_c_568_n 0.00353823f $X=4.81 $Y=1.765 $X2=0
+ $Y2=0
cc_327 N_A_27_368#_c_413_n N_VPWR_c_568_n 0.003573f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_328 N_A_27_368#_c_416_n N_VPWR_c_568_n 0.0102675f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_329 N_A_27_368#_c_417_n N_VPWR_c_568_n 0.033404f $X=1.46 $Y=2.475 $X2=0 $Y2=0
cc_330 N_A_27_368#_c_419_n N_A_348_368#_M1000_d 0.00826493f $X=2.36 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_331 N_A_27_368#_c_419_n N_A_348_368#_c_652_n 0.0281219f $X=2.36 $Y=2.145
+ $X2=0 $Y2=0
cc_332 N_A_27_368#_c_421_n N_A_348_368#_c_642_n 0.0134529f $X=2.445 $Y=2.06
+ $X2=0 $Y2=0
cc_333 N_A_27_368#_c_408_n N_A_348_368#_c_642_n 0.0137147f $X=3.82 $Y=1.485
+ $X2=0 $Y2=0
cc_334 N_A_27_368#_c_419_n N_A_348_368#_c_658_n 0.0133617f $X=2.36 $Y=2.145
+ $X2=0 $Y2=0
cc_335 N_A_27_368#_c_421_n N_A_348_368#_c_658_n 0.00484408f $X=2.445 $Y=2.06
+ $X2=0 $Y2=0
cc_336 N_A_27_368#_c_408_n N_A_348_368#_c_644_n 0.0452479f $X=3.82 $Y=1.485
+ $X2=0 $Y2=0
cc_337 N_A_27_368#_c_410_n N_A_348_368#_c_645_n 8.29946e-19 $X=3.91 $Y=1.765
+ $X2=0 $Y2=0
cc_338 N_A_27_368#_c_408_n N_A_348_368#_c_645_n 0.0209339f $X=3.82 $Y=1.485
+ $X2=0 $Y2=0
cc_339 N_A_27_368#_c_410_n N_A_348_368#_c_669_n 0.00637485f $X=3.91 $Y=1.765
+ $X2=0 $Y2=0
cc_340 N_A_27_368#_c_410_n N_A_348_368#_c_646_n 0.0128006f $X=3.91 $Y=1.765
+ $X2=0 $Y2=0
cc_341 N_A_27_368#_c_411_n N_A_348_368#_c_646_n 0.0128349f $X=4.36 $Y=1.765
+ $X2=0 $Y2=0
cc_342 N_A_27_368#_c_412_n N_A_348_368#_c_648_n 0.0128349f $X=4.81 $Y=1.765
+ $X2=0 $Y2=0
cc_343 N_A_27_368#_c_413_n N_A_348_368#_c_648_n 0.0135517f $X=5.26 $Y=1.765
+ $X2=0 $Y2=0
cc_344 N_A_27_368#_c_413_n N_A_348_368#_c_649_n 0.00799735f $X=5.26 $Y=1.765
+ $X2=0 $Y2=0
cc_345 N_A_27_368#_c_417_n N_A_348_368#_c_672_n 0.0133003f $X=1.46 $Y=2.475
+ $X2=0 $Y2=0
cc_346 N_A_27_368#_c_419_n N_A_348_368#_c_672_n 0.0131482f $X=2.36 $Y=2.145
+ $X2=0 $Y2=0
cc_347 N_A_27_368#_c_410_n N_Z_c_730_n 0.00218878f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_348 N_A_27_368#_c_411_n N_Z_c_730_n 6.83942e-19 $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_349 N_A_27_368#_c_405_n N_Z_c_730_n 0.0276567f $X=3.985 $Y=1.485 $X2=0 $Y2=0
cc_350 N_A_27_368#_c_409_n N_Z_c_730_n 0.00789892f $X=5.26 $Y=1.542 $X2=0 $Y2=0
cc_351 N_A_27_368#_c_410_n N_Z_c_734_n 0.00773563f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_352 N_A_27_368#_c_411_n N_Z_c_734_n 0.0085809f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_353 N_A_27_368#_c_412_n N_Z_c_734_n 5.86053e-19 $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_354 N_A_27_368#_M1005_g N_Z_c_742_n 0.00466922f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A_27_368#_M1013_g N_Z_c_742_n 0.00587139f $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_356 N_A_27_368#_M1014_g N_Z_c_742_n 5.63827e-19 $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A_27_368#_c_411_n N_Z_c_731_n 0.0120074f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_358 N_A_27_368#_c_412_n N_Z_c_731_n 0.0125823f $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_359 N_A_27_368#_c_518_p N_Z_c_731_n 0.0389377f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_360 N_A_27_368#_c_409_n N_Z_c_731_n 0.00762857f $X=5.26 $Y=1.542 $X2=0 $Y2=0
cc_361 N_A_27_368#_M1013_g N_Z_c_726_n 0.00891372f $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_362 N_A_27_368#_M1014_g N_Z_c_726_n 0.00944863f $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A_27_368#_c_518_p N_Z_c_726_n 0.0356525f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_364 N_A_27_368#_c_409_n N_Z_c_726_n 0.00224206f $X=5.26 $Y=1.542 $X2=0 $Y2=0
cc_365 N_A_27_368#_M1005_g N_Z_c_727_n 0.00373071f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A_27_368#_M1013_g N_Z_c_727_n 0.00235421f $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A_27_368#_c_518_p N_Z_c_727_n 0.0271537f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_368 N_A_27_368#_c_409_n N_Z_c_727_n 0.002312f $X=5.26 $Y=1.542 $X2=0 $Y2=0
cc_369 N_A_27_368#_M1013_g N_Z_c_757_n 5.63827e-19 $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A_27_368#_M1014_g N_Z_c_757_n 0.00640291f $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A_27_368#_M1019_g N_Z_c_757_n 0.0047509f $X=5.275 $Y=0.74 $X2=0 $Y2=0
cc_372 N_A_27_368#_M1014_g N_Z_c_728_n 0.00261386f $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A_27_368#_c_413_n N_Z_c_728_n 0.00291507f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_374 N_A_27_368#_M1019_g N_Z_c_728_n 0.00843462f $X=5.275 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A_27_368#_c_518_p N_Z_c_728_n 0.0214916f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_376 N_A_27_368#_c_409_n N_Z_c_728_n 0.0363865f $X=5.26 $Y=1.542 $X2=0 $Y2=0
cc_377 N_A_27_368#_M1014_g N_Z_c_729_n 0.00225227f $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A_27_368#_M1019_g N_Z_c_729_n 0.00363443f $X=5.275 $Y=0.74 $X2=0 $Y2=0
cc_379 N_A_27_368#_c_409_n N_Z_c_729_n 0.0013317f $X=5.26 $Y=1.542 $X2=0 $Y2=0
cc_380 N_A_27_368#_c_412_n Z 8.92358e-19 $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_381 N_A_27_368#_c_413_n Z 0.00211244f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_382 N_A_27_368#_c_409_n Z 0.00502298f $X=5.26 $Y=1.542 $X2=0 $Y2=0
cc_383 N_A_27_368#_c_411_n Z 5.85946e-19 $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_384 N_A_27_368#_c_412_n Z 0.0085809f $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_385 N_A_27_368#_c_413_n Z 0.00840931f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_386 N_A_27_368#_c_403_n N_VGND_c_794_n 0.024411f $X=0.32 $Y=0.515 $X2=0 $Y2=0
cc_387 N_A_27_368#_c_403_n N_VGND_c_801_n 0.0141895f $X=0.32 $Y=0.515 $X2=0
+ $Y2=0
cc_388 N_A_27_368#_M1005_g N_VGND_c_802_n 0.00278271f $X=3.965 $Y=0.74 $X2=0
+ $Y2=0
cc_389 N_A_27_368#_M1013_g N_VGND_c_802_n 0.00278271f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_390 N_A_27_368#_M1014_g N_VGND_c_802_n 0.00278271f $X=4.825 $Y=0.74 $X2=0
+ $Y2=0
cc_391 N_A_27_368#_M1019_g N_VGND_c_802_n 0.00278271f $X=5.275 $Y=0.74 $X2=0
+ $Y2=0
cc_392 N_A_27_368#_M1005_g N_VGND_c_803_n 0.00353526f $X=3.965 $Y=0.74 $X2=0
+ $Y2=0
cc_393 N_A_27_368#_M1013_g N_VGND_c_803_n 0.00353428f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_394 N_A_27_368#_M1014_g N_VGND_c_803_n 0.00353626f $X=4.825 $Y=0.74 $X2=0
+ $Y2=0
cc_395 N_A_27_368#_M1019_g N_VGND_c_803_n 0.00353613f $X=5.275 $Y=0.74 $X2=0
+ $Y2=0
cc_396 N_A_27_368#_c_403_n N_VGND_c_803_n 0.0117448f $X=0.32 $Y=0.515 $X2=0
+ $Y2=0
cc_397 N_A_27_368#_c_404_n N_A_378_74#_c_867_n 0.0137157f $X=2.53 $Y=1.565 $X2=0
+ $Y2=0
cc_398 N_A_27_368#_c_408_n N_A_378_74#_c_867_n 0.0195631f $X=3.82 $Y=1.485 $X2=0
+ $Y2=0
cc_399 N_A_27_368#_M1005_g N_A_378_74#_c_870_n 3.2654e-19 $X=3.965 $Y=0.74 $X2=0
+ $Y2=0
cc_400 N_A_27_368#_c_405_n N_A_378_74#_c_870_n 0.001265f $X=3.985 $Y=1.485 $X2=0
+ $Y2=0
cc_401 N_A_27_368#_c_408_n N_A_378_74#_c_870_n 0.0402638f $X=3.82 $Y=1.485 $X2=0
+ $Y2=0
cc_402 N_A_27_368#_c_409_n N_A_378_74#_c_870_n 3.70873e-19 $X=5.26 $Y=1.542
+ $X2=0 $Y2=0
cc_403 N_A_27_368#_M1005_g N_A_378_74#_c_871_n 0.0122971f $X=3.965 $Y=0.74 $X2=0
+ $Y2=0
cc_404 N_A_27_368#_M1013_g N_A_378_74#_c_871_n 0.0102404f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_405 N_A_27_368#_M1014_g N_A_378_74#_c_873_n 0.0103604f $X=4.825 $Y=0.74 $X2=0
+ $Y2=0
cc_406 N_A_27_368#_M1019_g N_A_378_74#_c_873_n 0.0139388f $X=5.275 $Y=0.74 $X2=0
+ $Y2=0
cc_407 N_A_27_368#_M1019_g N_A_378_74#_c_874_n 0.00159899f $X=5.275 $Y=0.74
+ $X2=0 $Y2=0
cc_408 N_A_27_368#_c_408_n N_A_378_74#_c_875_n 0.0134254f $X=3.82 $Y=1.485 $X2=0
+ $Y2=0
cc_409 N_VPWR_M1000_s N_A_348_368#_c_652_n 0.0037687f $X=2.185 $Y=1.84 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_570_n N_A_348_368#_c_652_n 0.0166605f $X=2.335 $Y=2.825 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_571_n N_A_348_368#_c_652_n 0.00216873f $X=3.07 $Y=3.33 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_573_n N_A_348_368#_c_652_n 0.00217512f $X=2.17 $Y=3.33 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_568_n N_A_348_368#_c_652_n 0.010241f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_414 N_VPWR_c_572_n N_A_348_368#_c_658_n 0.0152713f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_570_n N_A_348_368#_c_643_n 0.0156602f $X=2.335 $Y=2.825 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_571_n N_A_348_368#_c_643_n 0.00749631f $X=3.07 $Y=3.33 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_572_n N_A_348_368#_c_643_n 0.0261386f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_568_n N_A_348_368#_c_643_n 0.0062048f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_419 N_VPWR_M1002_s N_A_348_368#_c_644_n 0.00222494f $X=3.085 $Y=1.84 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_572_n N_A_348_368#_c_644_n 0.0154248f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_572_n N_A_348_368#_c_669_n 0.0488992f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_576_n N_A_348_368#_c_646_n 0.0441612f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_568_n N_A_348_368#_c_646_n 0.0249452f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_572_n N_A_348_368#_c_647_n 0.012272f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_576_n N_A_348_368#_c_647_n 0.017869f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_426 N_VPWR_c_568_n N_A_348_368#_c_647_n 0.00965079f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_576_n N_A_348_368#_c_648_n 0.0620829f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_568_n N_A_348_368#_c_648_n 0.0346647f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_570_n N_A_348_368#_c_672_n 0.00521095f $X=2.335 $Y=2.825 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_573_n N_A_348_368#_c_672_n 0.00421509f $X=2.17 $Y=3.33 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_568_n N_A_348_368#_c_672_n 0.00547139f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_572_n N_A_348_368#_c_713_n 0.0121475f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_576_n N_A_348_368#_c_650_n 0.016488f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_568_n N_A_348_368#_c_650_n 0.00894187f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_435 N_A_348_368#_c_646_n N_Z_M1004_d 0.00197722f $X=4.47 $Y=2.99 $X2=0 $Y2=0
cc_436 N_A_348_368#_c_648_n N_Z_M1010_d 0.00197722f $X=5.4 $Y=2.99 $X2=0 $Y2=0
cc_437 N_A_348_368#_c_645_n N_Z_c_730_n 0.013128f $X=3.645 $Y=1.99 $X2=0 $Y2=0
cc_438 N_A_348_368#_c_669_n N_Z_c_734_n 0.049886f $X=3.685 $Y=2.815 $X2=0 $Y2=0
cc_439 N_A_348_368#_c_646_n N_Z_c_734_n 0.0160777f $X=4.47 $Y=2.99 $X2=0 $Y2=0
cc_440 N_A_348_368#_M1008_s N_Z_c_731_n 0.00197722f $X=4.435 $Y=1.84 $X2=0 $Y2=0
cc_441 N_A_348_368#_c_722_p N_Z_c_731_n 0.0151327f $X=4.585 $Y=2.325 $X2=0 $Y2=0
cc_442 N_A_348_368#_c_649_n Z 0.0123713f $X=5.485 $Y=1.985 $X2=0 $Y2=0
cc_443 N_A_348_368#_c_648_n Z 0.0164339f $X=5.4 $Y=2.99 $X2=0 $Y2=0
cc_444 N_A_348_368#_c_649_n Z 0.0509581f $X=5.485 $Y=1.985 $X2=0 $Y2=0
cc_445 N_Z_c_726_n N_A_378_74#_M1013_d 0.00176461f $X=4.875 $Y=1.065 $X2=0 $Y2=0
cc_446 N_Z_c_727_n N_A_378_74#_c_870_n 0.00862188f $X=4.345 $Y=1.065 $X2=0 $Y2=0
cc_447 N_Z_M1005_s N_A_378_74#_c_871_n 0.00176461f $X=4.04 $Y=0.37 $X2=0 $Y2=0
cc_448 N_Z_c_742_n N_A_378_74#_c_871_n 0.0158052f $X=4.18 $Y=0.82 $X2=0 $Y2=0
cc_449 N_Z_c_726_n N_A_378_74#_c_871_n 0.0031794f $X=4.875 $Y=1.065 $X2=0 $Y2=0
cc_450 N_Z_c_726_n N_A_378_74#_c_923_n 0.0132844f $X=4.875 $Y=1.065 $X2=0 $Y2=0
cc_451 N_Z_M1014_s N_A_378_74#_c_873_n 0.00197722f $X=4.9 $Y=0.37 $X2=0 $Y2=0
cc_452 N_Z_c_726_n N_A_378_74#_c_873_n 0.0031794f $X=4.875 $Y=1.065 $X2=0 $Y2=0
cc_453 N_Z_c_757_n N_A_378_74#_c_873_n 0.0160331f $X=5.04 $Y=0.86 $X2=0 $Y2=0
cc_454 N_Z_c_729_n N_A_378_74#_c_874_n 0.00622221f $X=5.04 $Y=1.065 $X2=0 $Y2=0
cc_455 N_VGND_c_795_n N_A_378_74#_c_866_n 0.0229082f $X=2.46 $Y=0.515 $X2=0
+ $Y2=0
cc_456 N_VGND_c_797_n N_A_378_74#_c_866_n 0.00749631f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_457 N_VGND_c_803_n N_A_378_74#_c_866_n 0.0062048f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_458 N_VGND_c_795_n N_A_378_74#_c_867_n 0.0216086f $X=2.46 $Y=0.515 $X2=0
+ $Y2=0
cc_459 N_VGND_c_795_n N_A_378_74#_c_869_n 0.0229082f $X=2.46 $Y=0.515 $X2=0
+ $Y2=0
cc_460 N_VGND_c_796_n N_A_378_74#_c_869_n 0.0164868f $X=3.32 $Y=0.645 $X2=0
+ $Y2=0
cc_461 N_VGND_c_799_n N_A_378_74#_c_869_n 0.00749631f $X=3.155 $Y=0 $X2=0 $Y2=0
cc_462 N_VGND_c_803_n N_A_378_74#_c_869_n 0.0062048f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_M1009_d N_A_378_74#_c_870_n 0.00176461f $X=3.18 $Y=0.37 $X2=0
+ $Y2=0
cc_464 N_VGND_c_796_n N_A_378_74#_c_870_n 0.0152916f $X=3.32 $Y=0.645 $X2=0
+ $Y2=0
cc_465 N_VGND_c_802_n N_A_378_74#_c_871_n 0.043517f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_466 N_VGND_c_803_n N_A_378_74#_c_871_n 0.0245693f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_467 N_VGND_c_796_n N_A_378_74#_c_872_n 0.0112234f $X=3.32 $Y=0.645 $X2=0
+ $Y2=0
cc_468 N_VGND_c_802_n N_A_378_74#_c_872_n 0.0178338f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_803_n N_A_378_74#_c_872_n 0.00960503f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_c_802_n N_A_378_74#_c_873_n 0.0627271f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_803_n N_A_378_74#_c_873_n 0.0350406f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_c_802_n N_A_378_74#_c_876_n 0.0120038f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_803_n N_A_378_74#_c_876_n 0.00657483f $X=5.52 $Y=0 $X2=0 $Y2=0
