# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dlxbn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dlxbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.260000 0.835000 1.930000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.765000 1.820000 6.130000 2.980000 ;
        RECT 5.790000 0.350000 6.130000 1.100000 ;
        RECT 5.960000 1.100000 6.130000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.537600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715000 0.350000 8.050000 2.980000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.690000 1.335000 2.150000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 0.410000 ;
        RECT 2.340000  0.085000 2.675000 0.410000 ;
        RECT 4.705000  0.085000 5.035000 0.960000 ;
        RECT 6.300000  0.085000 6.550000 1.130000 ;
        RECT 7.290000  0.085000 7.540000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.735000 2.320000 1.065000 3.245000 ;
        RECT 2.380000 2.730000 2.710000 3.245000 ;
        RECT 4.480000 2.060000 5.020000 3.245000 ;
        RECT 6.300000 2.100000 6.550000 3.245000 ;
        RECT 7.265000 1.820000 7.515000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.580000 2.865000 0.750000 ;
      RECT 0.095000 0.750000 0.445000 1.090000 ;
      RECT 0.095000 1.090000 0.265000 2.100000 ;
      RECT 0.095000 2.100000 0.545000 2.980000 ;
      RECT 1.135000 0.920000 1.465000 1.260000 ;
      RECT 1.135000 1.260000 1.905000 1.520000 ;
      RECT 1.235000 2.320000 1.675000 2.390000 ;
      RECT 1.235000 2.390000 4.145000 2.560000 ;
      RECT 1.235000 2.560000 1.565000 2.980000 ;
      RECT 1.505000 1.520000 1.675000 2.320000 ;
      RECT 1.695000 0.920000 2.245000 1.090000 ;
      RECT 1.845000 1.880000 2.910000 2.220000 ;
      RECT 2.075000 1.090000 2.245000 1.710000 ;
      RECT 2.075000 1.710000 3.340000 1.880000 ;
      RECT 2.535000 0.750000 2.865000 1.510000 ;
      RECT 3.035000 0.255000 4.260000 0.505000 ;
      RECT 3.035000 0.505000 3.205000 1.470000 ;
      RECT 3.035000 1.470000 3.340000 1.710000 ;
      RECT 3.260000 2.050000 3.805000 2.220000 ;
      RECT 3.375000 0.725000 4.135000 1.055000 ;
      RECT 3.510000 1.055000 4.135000 1.130000 ;
      RECT 3.510000 1.130000 5.220000 1.300000 ;
      RECT 3.510000 1.300000 3.680000 2.050000 ;
      RECT 3.850000 1.470000 4.145000 1.800000 ;
      RECT 3.975000 1.800000 4.145000 2.390000 ;
      RECT 4.315000 1.470000 4.645000 1.720000 ;
      RECT 4.315000 1.720000 5.560000 1.890000 ;
      RECT 4.890000 1.300000 5.220000 1.550000 ;
      RECT 5.205000 0.350000 5.560000 0.960000 ;
      RECT 5.220000 1.890000 5.560000 2.900000 ;
      RECT 5.390000 0.960000 5.560000 1.270000 ;
      RECT 5.390000 1.270000 5.790000 1.600000 ;
      RECT 5.390000 1.600000 5.560000 1.720000 ;
      RECT 6.720000 0.540000 7.060000 1.300000 ;
      RECT 6.720000 1.300000 7.500000 1.630000 ;
      RECT 6.720000 1.630000 7.065000 2.980000 ;
  END
END sky130_fd_sc_hs__dlxbn_1
