* NGSPICE file created from sky130_fd_sc_hs__mux2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux2_2 A0 A1 S VGND VNB VPB VPWR X
M1000 X a_116_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=1.2092e+12p ps=8.77e+06u
M1001 VPWR a_116_368# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR S a_459_48# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1003 a_116_368# A0 a_38_74# VNB nlowvt w=740000u l=150000u
+  ad=4.255e+11p pd=2.63e+06u as=4.292e+11p ps=4.12e+06u
M1004 X a_116_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=9.4915e+11p ps=7.09e+06u
M1005 a_38_74# a_459_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_270_74# A1 a_116_368# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1007 a_206_368# A1 a_116_368# VPB pshort w=1e+06u l=150000u
+  ad=5.9e+11p pd=5.18e+06u as=3e+11p ps=2.6e+06u
M1008 a_116_368# A0 a_27_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=5.9e+11p ps=5.18e+06u
M1009 a_206_368# a_459_48# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND S a_270_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR S a_27_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND S a_459_48# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 VGND a_116_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

