* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux2_4 A0 A1 S VGND VNB VPB VPWR X
X0 a_27_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_722_391# A0 a_193_241# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_722_391# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X3 VGND a_27_368# a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_193_241# A1 a_936_391# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_709_119# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_709_119# A1 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 VPWR a_27_368# a_936_391# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_193_241# A0 a_722_391# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X12 a_937_119# A0 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_936_391# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X14 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 VPWR S a_722_391# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X17 a_936_391# A1 a_193_241# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X18 a_193_241# A0 a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_193_241# A1 a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X21 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_27_368# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 a_937_119# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X25 VGND S a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
