* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_509_392# S1 a_2199_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_2199_74# a_2489_347# a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_116_392# a_758_306# a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X3 a_1285_377# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 a_1450_121# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_1278_121# a_758_306# a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_1285_377# a_758_306# a_1191_121# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 VGND A2 a_1278_121# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_1465_377# S0 a_1191_121# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X9 a_2199_74# a_2489_347# a_1191_121# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 VPWR A2 a_1465_377# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X11 a_509_392# a_2489_347# a_2199_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_509_392# a_758_306# a_299_126# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_758_306# S0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X14 a_114_126# S0 a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 VPWR A1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X16 a_296_392# S0 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X17 a_509_392# S0 a_114_126# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 a_1450_121# S0 a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 VGND A3 a_1450_121# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_1191_121# S0 a_1450_121# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 a_1191_121# a_2489_347# a_2199_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X22 VPWR a_2199_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X23 a_1278_121# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 a_758_306# S0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_2199_74# S1 a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X26 VPWR A0 a_296_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X27 a_509_392# a_758_306# a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X28 VGND A1 a_114_126# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X29 X a_2199_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X30 X a_2199_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 VGND A0 a_299_126# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X32 a_299_126# a_758_306# a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X33 a_2489_347# S1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 a_1191_121# a_758_306# a_1285_377# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X35 a_1191_121# S1 a_2199_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X36 a_114_126# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X37 X a_2199_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 a_1191_121# S0 a_1465_377# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X39 a_296_392# A0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X40 a_509_392# S0 a_296_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X41 VPWR A3 a_1285_377# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X42 X a_2199_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X43 VGND a_2199_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X44 VGND a_2199_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X45 a_1465_377# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X46 a_2199_74# S1 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X47 a_299_126# A0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X48 a_2489_347# S1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X49 a_1191_121# a_758_306# a_1278_121# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X50 a_116_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X51 VPWR a_2199_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
.ends
