* File: sky130_fd_sc_hs__dlrbn_1.pex.spice
* Created: Tue Sep  1 20:01:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DLRBN_1%D 2 5 7 9 10 13
r33 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.425
+ $X2=0.59 $Y2=1.26
r34 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6
+ $Y=1.425 $X2=0.6 $Y2=1.425
r35 10 14 2.24265 $w=6.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.58 $X2=0.6
+ $Y2=1.58
r36 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
r37 5 15 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.5 $Y=0.835 $X2=0.5
+ $Y2=1.26
r38 2 7 49.5674 $w=2.82e-07 $l=3.29773e-07 $layer=POLY_cond $X=0.59 $Y=1.755
+ $X2=0.505 $Y2=2.045
r39 1 13 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.59 $Y=1.435 $X2=0.59
+ $Y2=1.425
r40 1 2 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.59 $Y=1.435 $X2=0.59
+ $Y2=1.755
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%GATE_N 3 6 7 9 10 13 14
r35 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.425
+ $X2=1.18 $Y2=1.26
r36 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.425 $X2=1.17 $Y2=1.425
r37 10 14 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.425
r38 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.265 $Y=2.045
+ $X2=1.265 $Y2=2.54
r39 6 7 49.5674 $w=2.82e-07 $l=3.29773e-07 $layer=POLY_cond $X=1.18 $Y=1.755
+ $X2=1.265 $Y2=2.045
r40 5 13 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=1.18 $Y=1.435 $X2=1.18
+ $Y2=1.425
r41 5 6 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.18 $Y=1.435 $X2=1.18
+ $Y2=1.755
r42 3 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.08 $Y=0.74 $X2=1.08
+ $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%A_231_74# 1 2 9 11 12 14 17 18 20 23 26 27
+ 30 32 33 34 37 41 44 45 49 53 57 59 63 66 69 71
c160 53 0 9.3463e-20 $X=2.35 $Y=1.385
c161 26 0 5.58535e-20 $X=2.47 $Y=2.22
r162 63 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.445 $Y=1.285
+ $X2=3.445 $Y2=1.12
r163 62 64 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=1.285
+ $X2=3.445 $Y2=1.45
r164 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.285 $X2=3.445 $Y2=1.285
r165 59 62 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=3.445 $Y=1.215
+ $X2=3.445 $Y2=1.285
r166 55 57 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.205 $Y=2.055
+ $X2=3.365 $Y2=2.055
r167 53 67 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.332 $Y=1.385
+ $X2=2.332 $Y2=1.55
r168 53 66 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.332 $Y=1.385
+ $X2=2.332 $Y2=1.22
r169 52 54 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=1.385
+ $X2=2.37 $Y2=1.55
r170 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.35
+ $Y=1.385 $X2=2.35 $Y2=1.385
r171 49 52 5.29501 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.37 $Y=1.215
+ $X2=2.37 $Y2=1.385
r172 44 47 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.54 $Y=2.305
+ $X2=1.54 $Y2=2.33
r173 44 45 10.3232 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.54 $Y=2.305
+ $X2=1.54 $Y2=2.1
r174 43 45 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.59 $Y=1.09
+ $X2=1.59 $Y2=2.1
r175 41 43 18.7979 $w=5.43e-07 $l=5.75e-07 $layer=LI1_cond $X=1.402 $Y=0.515
+ $X2=1.402 $Y2=1.09
r176 38 71 25.1593 $w=3.64e-07 $l=1.9e-07 $layer=POLY_cond $X=4.125 $Y=2.257
+ $X2=3.935 $Y2=2.257
r177 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.125
+ $Y=2.215 $X2=4.125 $Y2=2.215
r178 35 37 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=4.125 $Y=2.905
+ $X2=4.125 $Y2=2.215
r179 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.96 $Y=2.99
+ $X2=4.125 $Y2=2.905
r180 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.96 $Y=2.99
+ $X2=3.29 $Y2=2.99
r181 32 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=1.97
+ $X2=3.365 $Y2=2.055
r182 32 64 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.365 $Y=1.97
+ $X2=3.365 $Y2=1.45
r183 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.205 $Y=2.905
+ $X2=3.29 $Y2=2.99
r184 29 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=2.14
+ $X2=3.205 $Y2=2.055
r185 29 30 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.205 $Y=2.14
+ $X2=3.205 $Y2=2.905
r186 28 49 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.555 $Y=1.215
+ $X2=2.37 $Y2=1.215
r187 27 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=1.215
+ $X2=3.445 $Y2=1.215
r188 27 28 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.28 $Y=1.215
+ $X2=2.555 $Y2=1.215
r189 26 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.47 $Y=2.22
+ $X2=2.47 $Y2=1.55
r190 24 44 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.675 $Y=2.305
+ $X2=1.54 $Y2=2.305
r191 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.385 $Y=2.305
+ $X2=2.47 $Y2=2.22
r192 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.385 $Y=2.305
+ $X2=1.675 $Y2=2.305
r193 18 71 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.935 $Y=2.465
+ $X2=3.935 $Y2=2.257
r194 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.935 $Y=2.465
+ $X2=3.935 $Y2=2.75
r195 17 69 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.355 $Y=0.69
+ $X2=3.355 $Y2=1.12
r196 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.36 $Y=1.885
+ $X2=2.36 $Y2=2.38
r197 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.36 $Y=1.795
+ $X2=2.36 $Y2=1.885
r198 11 67 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=2.36 $Y=1.795
+ $X2=2.36 $Y2=1.55
r199 9 66 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.225 $Y=0.74
+ $X2=2.225 $Y2=1.22
r200 2 47 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.12 $X2=1.49 $Y2=2.33
r201 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.37 $X2=1.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%A_27_424# 1 2 9 11 13 14 18 21 23 26 27 28
+ 29 32 33 34 35 40
c108 40 0 2.24964e-19 $X=2.905 $Y=1.635
c109 32 0 8.30347e-20 $X=2.825 $Y=2.56
r110 40 43 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=1.635
+ $X2=2.905 $Y2=1.8
r111 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=1.635 $X2=2.905 $Y2=1.635
r112 35 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.93 $Y=2.645
+ $X2=1.93 $Y2=2.815
r113 32 43 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.825 $Y=2.56
+ $X2=2.825 $Y2=1.8
r114 30 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=2.645
+ $X2=1.93 $Y2=2.645
r115 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.74 $Y=2.645
+ $X2=2.825 $Y2=2.56
r116 29 30 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.74 $Y=2.645
+ $X2=2.015 $Y2=2.645
r117 27 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=2.815
+ $X2=1.93 $Y2=2.815
r118 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.845 $Y=2.815
+ $X2=1.235 $Y2=2.815
r119 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.73
+ $X2=1.235 $Y2=2.815
r120 25 26 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.15 $Y=2.24
+ $X2=1.15 $Y2=2.73
r121 24 34 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.365 $Y=2.155
+ $X2=0.23 $Y2=2.155
r122 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=2.155
+ $X2=1.15 $Y2=2.24
r123 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.065 $Y=2.155
+ $X2=0.365 $Y2=2.155
r124 19 34 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=2.24
+ $X2=0.23 $Y2=2.155
r125 19 21 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.23 $Y=2.24
+ $X2=0.23 $Y2=2.265
r126 18 34 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.18 $Y=2.07
+ $X2=0.23 $Y2=2.155
r127 18 33 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.18 $Y=2.07
+ $X2=0.18 $Y2=1.09
r128 14 33 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=0.272 $Y=0.913
+ $X2=0.272 $Y2=1.09
r129 14 16 3.36789 $w=3.55e-07 $l=9.8e-08 $layer=LI1_cond $X=0.272 $Y=0.913
+ $X2=0.272 $Y2=0.815
r130 11 41 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.98 $Y=1.885
+ $X2=2.905 $Y2=1.635
r131 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.98 $Y=1.885
+ $X2=2.98 $Y2=2.46
r132 7 41 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.965 $Y=1.47
+ $X2=2.905 $Y2=1.635
r133 7 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.965 $Y=1.47
+ $X2=2.965 $Y2=0.69
r134 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r135 1 16 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.56 $X2=0.285 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%A_373_74# 1 2 7 9 10 11 13 16 19 22 23 27 28
+ 30 34 37
c99 23 0 1.8903e-19 $X=3.875 $Y=0.865
c100 11 0 2.14535e-19 $X=3.49 $Y=1.765
r101 31 34 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.93 $Y=1.885
+ $X2=2.05 $Y2=1.885
r102 28 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.04 $Y=1.285
+ $X2=4.04 $Y2=1.45
r103 28 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.04 $Y=1.285
+ $X2=4.04 $Y2=1.12
r104 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.04
+ $Y=1.285 $X2=4.04 $Y2=1.285
r105 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.04 $Y=0.95
+ $X2=4.04 $Y2=1.285
r106 24 30 2.76166 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.175 $Y=0.865
+ $X2=2.01 $Y2=0.87
r107 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=0.865
+ $X2=4.04 $Y2=0.95
r108 23 24 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=3.875 $Y=0.865
+ $X2=2.175 $Y2=0.865
r109 22 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=1.72
+ $X2=1.93 $Y2=1.885
r110 21 30 3.70735 $w=2.5e-07 $l=1.23693e-07 $layer=LI1_cond $X=1.93 $Y=0.96
+ $X2=2.01 $Y2=0.87
r111 21 22 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.93 $Y=0.96
+ $X2=1.93 $Y2=1.72
r112 17 30 3.70735 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.01 $Y=0.78 $X2=2.01
+ $Y2=0.87
r113 17 19 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.01 $Y=0.78
+ $X2=2.01 $Y2=0.515
r114 16 37 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.13 $Y=0.8
+ $X2=4.13 $Y2=1.12
r115 13 38 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.95 $Y=1.69
+ $X2=3.95 $Y2=1.45
r116 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.95 $Y2=1.69
r117 10 11 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.49 $Y2=1.765
r118 7 11 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=3.4 $Y=1.885
+ $X2=3.49 $Y2=1.765
r119 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.4 $Y=1.885 $X2=3.4
+ $Y2=2.46
r120 2 34 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.74 $X2=2.05 $Y2=1.885
r121 1 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.865
+ $Y=0.37 $X2=2.01 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%A_889_92# 1 2 9 11 13 14 16 17 19 20 22 23
+ 25 27 29 37 40 43 45 48 49 51 54 58
c128 48 0 1.12758e-19 $X=6.435 $Y=1.72
c129 17 0 1.37399e-19 $X=6.535 $Y=1.635
c130 9 0 1.8903e-19 $X=4.52 $Y=0.8
r131 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.645
+ $Y=1.385 $X2=6.645 $Y2=1.385
r132 55 58 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.435 $Y=1.385
+ $X2=6.645 $Y2=1.385
r133 53 54 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.78 $Y=2.005
+ $X2=5.945 $Y2=2.005
r134 50 53 8.49845 $w=5.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.375 $Y=2.005
+ $X2=5.78 $Y2=2.005
r135 50 51 3.88629 $w=5.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=2.005
+ $X2=5.29 $Y2=2.005
r136 47 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=1.55
+ $X2=6.435 $Y2=1.385
r137 47 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.435 $Y=1.55
+ $X2=6.435 $Y2=1.72
r138 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.35 $Y=1.805
+ $X2=6.435 $Y2=1.72
r139 45 54 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.35 $Y=1.805
+ $X2=5.945 $Y2=1.805
r140 41 53 3.93508 $w=3.3e-07 $l=2.85e-07 $layer=LI1_cond $X=5.78 $Y=2.29
+ $X2=5.78 $Y2=2.005
r141 41 43 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=5.78 $Y=2.29
+ $X2=5.78 $Y2=2.685
r142 40 50 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=5.375 $Y=1.72
+ $X2=5.375 $Y2=2.005
r143 40 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.375 $Y=1.72
+ $X2=5.375 $Y2=1.05
r144 35 49 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.335 $Y=0.925
+ $X2=5.335 $Y2=1.05
r145 35 37 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=5.335 $Y=0.925
+ $X2=5.335 $Y2=0.515
r146 32 51 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=4.695 $Y=2.125
+ $X2=5.29 $Y2=2.125
r147 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.695
+ $Y=2.125 $X2=4.695 $Y2=2.125
r148 29 59 100.982 $w=3.6e-07 $l=6.3e-07 $layer=POLY_cond $X=7.275 $Y=1.4
+ $X2=6.645 $Y2=1.4
r149 28 29 3.99919 $w=3.6e-07 $l=2.05e-07 $layer=POLY_cond $X=7.48 $Y=1.4
+ $X2=7.275 $Y2=1.4
r150 26 59 3.20579 $w=3.6e-07 $l=2e-08 $layer=POLY_cond $X=6.625 $Y=1.4
+ $X2=6.645 $Y2=1.4
r151 26 27 6.023 $w=3.6e-07 $l=1.02616e-07 $layer=POLY_cond $X=6.625 $Y=1.4
+ $X2=6.535 $Y2=1.427
r152 23 28 41.0971 $w=3.78e-07 $l=2.3622e-07 $layer=POLY_cond $X=7.61 $Y=1.22
+ $X2=7.48 $Y2=1.4
r153 23 25 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.61 $Y=1.22
+ $X2=7.61 $Y2=0.835
r154 20 28 74.8881 $w=3.78e-07 $l=4.99199e-07 $layer=POLY_cond $X=7.595 $Y=1.845
+ $X2=7.48 $Y2=1.4
r155 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.595 $Y=1.845
+ $X2=7.595 $Y2=2.34
r156 17 27 39.2672 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.535 $Y=1.635
+ $X2=6.535 $Y2=1.427
r157 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.535 $Y=1.635
+ $X2=6.535 $Y2=2.27
r158 14 27 39.2672 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=6.52 $Y=1.22
+ $X2=6.535 $Y2=1.427
r159 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.52 $Y=1.22
+ $X2=6.52 $Y2=0.74
r160 11 33 73.3766 $w=2.49e-07 $l=3.5564e-07 $layer=POLY_cond $X=4.62 $Y=2.465
+ $X2=4.652 $Y2=2.125
r161 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.62 $Y=2.465
+ $X2=4.62 $Y2=2.75
r162 7 33 91.7662 $w=2.49e-07 $l=4.96634e-07 $layer=POLY_cond $X=4.52 $Y=1.69
+ $X2=4.652 $Y2=2.125
r163 7 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=4.52 $Y=1.69 $X2=4.52
+ $Y2=0.8
r164 2 53 400 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_PDIFF $count=1 $X=5.62
+ $Y=1.71 $X2=5.78 $Y2=1.885
r165 2 43 400 $w=1.7e-07 $l=1.05196e-06 $layer=licon1_PDIFF $count=1 $X=5.62
+ $Y=1.71 $X2=5.78 $Y2=2.685
r166 1 37 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.23
+ $Y=0.37 $X2=5.375 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%A_686_74# 1 2 7 9 10 12 14 15 21 22 27 31 32
+ 34 35
r93 34 36 10.5366 $w=3.48e-07 $l=3.2e-07 $layer=LI1_cond $X=4.55 $Y=1.385
+ $X2=4.55 $Y2=1.705
r94 34 35 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.55 $Y=1.385
+ $X2=4.55 $Y2=1.22
r95 31 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=2.57
+ $X2=3.625 $Y2=2.405
r96 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.005
+ $Y=1.385 $X2=5.005 $Y2=1.385
r97 25 34 1.07274 $w=3.3e-07 $l=1.75e-07 $layer=LI1_cond $X=4.725 $Y=1.385
+ $X2=4.55 $Y2=1.385
r98 25 27 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.725 $Y=1.385
+ $X2=5.005 $Y2=1.385
r99 23 35 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.46 $Y=0.61
+ $X2=4.46 $Y2=1.22
r100 21 36 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.375 $Y=1.705
+ $X2=4.55 $Y2=1.705
r101 21 22 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.375 $Y=1.705
+ $X2=3.79 $Y2=1.705
r102 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.705 $Y=1.79
+ $X2=3.79 $Y2=1.705
r103 19 32 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.705 $Y=1.79
+ $X2=3.705 $Y2=2.405
r104 15 23 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.375 $Y=0.485
+ $X2=4.46 $Y2=0.61
r105 15 17 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=4.375 $Y=0.485
+ $X2=3.72 $Y2=0.485
r106 14 28 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=5.455 $Y=1.385
+ $X2=5.005 $Y2=1.385
r107 10 14 44.1289 $w=1.9e-07 $l=1.79374e-07 $layer=POLY_cond $X=5.59 $Y=1.22
+ $X2=5.56 $Y2=1.385
r108 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.59 $Y=1.22
+ $X2=5.59 $Y2=0.74
r109 7 14 65.692 $w=1.9e-07 $l=2.57391e-07 $layer=POLY_cond $X=5.545 $Y=1.635
+ $X2=5.56 $Y2=1.385
r110 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.545 $Y=1.635
+ $X2=5.545 $Y2=2.27
r111 2 31 600 $w=1.7e-07 $l=6.80882e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.96 $X2=3.625 $Y2=2.57
r112 1 17 182 $w=1.7e-07 $l=3.59235e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.37 $X2=3.72 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%RESET_B 1 3 4 6 7
c31 1 0 1.84321e-19 $X=5.98 $Y=1.22
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.04
+ $Y=1.385 $X2=6.04 $Y2=1.385
r33 7 11 3.40065 $w=3.03e-07 $l=9e-08 $layer=LI1_cond $X=6.027 $Y=1.295
+ $X2=6.027 $Y2=1.385
r34 4 10 52.2586 $w=2.99e-07 $l=2.66927e-07 $layer=POLY_cond $X=6.005 $Y=1.635
+ $X2=6.04 $Y2=1.385
r35 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.005 $Y=1.635
+ $X2=6.005 $Y2=2.27
r36 1 10 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.98 $Y=1.22
+ $X2=6.04 $Y2=1.385
r37 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.98 $Y=1.22 $X2=5.98
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%A_1437_112# 1 2 9 11 13 16 20 24 27
c38 20 0 1.37399e-19 $X=7.37 $Y=2.065
r39 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.06
+ $Y=1.465 $X2=8.06 $Y2=1.465
r40 22 27 0.533013 $w=3.3e-07 $l=1.38e-07 $layer=LI1_cond $X=7.56 $Y=1.465
+ $X2=7.422 $Y2=1.465
r41 22 24 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=7.56 $Y=1.465 $X2=8.06
+ $Y2=1.465
r42 18 27 6.22203 $w=2.62e-07 $l=1.70895e-07 $layer=LI1_cond $X=7.41 $Y=1.63
+ $X2=7.422 $Y2=1.465
r43 18 20 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=7.41 $Y=1.63
+ $X2=7.41 $Y2=2.065
r44 14 27 6.22203 $w=2.62e-07 $l=1.65e-07 $layer=LI1_cond $X=7.422 $Y=1.3
+ $X2=7.422 $Y2=1.465
r45 14 16 19.4868 $w=2.73e-07 $l=4.65e-07 $layer=LI1_cond $X=7.422 $Y=1.3
+ $X2=7.422 $Y2=0.835
r46 11 25 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.06 $Y2=1.465
r47 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=2.4
r48 7 25 38.6549 $w=2.86e-07 $l=1.94808e-07 $layer=POLY_cond $X=8.125 $Y=1.3
+ $X2=8.06 $Y2=1.465
r49 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.125 $Y=1.3 $X2=8.125
+ $Y2=0.74
r50 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=7.245
+ $Y=1.92 $X2=7.37 $Y2=2.065
r51 1 16 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.56 $X2=7.395 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%VPWR 1 2 3 4 5 18 22 26 30 35 36 37 39 44 52
+ 64 73 74 77 80 83 90
c104 4 0 1.12758e-19 $X=6.08 $Y=1.71
r105 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 74 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r109 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r110 71 90 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.01 $Y=3.33
+ $X2=7.877 $Y2=3.33
r111 71 73 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.01 $Y=3.33
+ $X2=8.4 $Y2=3.33
r112 70 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r117 64 90 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.745 $Y=3.33
+ $X2=7.877 $Y2=3.33
r118 64 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=3.33
+ $X2=7.44 $Y2=3.33
r119 63 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r120 63 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r121 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r122 60 62 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.445 $Y=3.33
+ $X2=6 $Y2=3.33
r123 59 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r124 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 56 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r126 55 58 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r128 53 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.67 $Y2=3.33
r129 53 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.12 $Y2=3.33
r130 52 60 9.90988 $w=1.7e-07 $l=3.83e-07 $layer=LI1_cond $X=5.062 $Y=3.33
+ $X2=5.445 $Y2=3.33
r131 52 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r132 52 83 10.0846 $w=7.63e-07 $l=6.45e-07 $layer=LI1_cond $X=5.062 $Y=3.33
+ $X2=5.062 $Y2=2.685
r133 52 58 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.68 $Y=3.33
+ $X2=4.56 $Y2=3.33
r134 51 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r139 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 45 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r141 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 44 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.67 $Y2=3.33
r143 44 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r144 42 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r145 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 39 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r147 39 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r148 37 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r149 37 56 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=3.12 $Y2=3.33
r150 35 62 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.115 $Y=3.33
+ $X2=6 $Y2=3.33
r151 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=3.33
+ $X2=6.28 $Y2=3.33
r152 34 66 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.445 $Y=3.33
+ $X2=6.48 $Y2=3.33
r153 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=3.33
+ $X2=6.28 $Y2=3.33
r154 30 33 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=7.877 $Y=1.985
+ $X2=7.877 $Y2=2.815
r155 28 90 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.877 $Y=3.245
+ $X2=7.877 $Y2=3.33
r156 28 33 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=7.877 $Y=3.245
+ $X2=7.877 $Y2=2.815
r157 24 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=3.245
+ $X2=6.28 $Y2=3.33
r158 24 26 38.4148 $w=3.28e-07 $l=1.1e-06 $layer=LI1_cond $X=6.28 $Y=3.245
+ $X2=6.28 $Y2=2.145
r159 20 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=3.33
r160 20 22 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=2.985
r161 16 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r162 16 18 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.495
r163 5 33 600 $w=1.7e-07 $l=1.00788e-06 $layer=licon1_PDIFF $count=1 $X=7.67
+ $Y=1.92 $X2=7.91 $Y2=2.815
r164 5 30 300 $w=1.7e-07 $l=2.70555e-07 $layer=licon1_PDIFF $count=2 $X=7.67
+ $Y=1.92 $X2=7.91 $Y2=1.985
r165 4 26 300 $w=1.7e-07 $l=5.25571e-07 $layer=licon1_PDIFF $count=2 $X=6.08
+ $Y=1.71 $X2=6.28 $Y2=2.145
r166 3 83 300 $w=1.7e-07 $l=6.53491e-07 $layer=licon1_PDIFF $count=2 $X=4.695
+ $Y=2.54 $X2=5.28 $Y2=2.685
r167 2 22 600 $w=1.7e-07 $l=1.13644e-06 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.96 $X2=2.67 $Y2=2.985
r168 1 18 300 $w=1.7e-07 $l=4.43706e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.12 $X2=0.73 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%Q 1 2 11 12 13 14 15 16 29
c33 29 0 1.84321e-19 $X=6.735 $Y=0.515
r34 16 26 7.59257 $w=4.23e-07 $l=2.8e-07 $layer=LI1_cond $X=6.902 $Y=2.405
+ $X2=6.902 $Y2=2.685
r35 15 16 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=6.902 $Y=2.035
+ $X2=6.902 $Y2=2.405
r36 14 35 8.96211 $w=5.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.84 $Y=0.925
+ $X2=6.84 $Y2=1.05
r37 13 14 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=6.84 $Y=0.555
+ $X2=6.84 $Y2=0.925
r38 13 29 0.869875 $w=5.48e-07 $l=4e-08 $layer=LI1_cond $X=6.84 $Y=0.555
+ $X2=6.84 $Y2=0.515
r39 12 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.03 $Y=1.72
+ $X2=7.03 $Y2=1.05
r40 11 12 8.76046 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=6.902 $Y=1.885
+ $X2=6.902 $Y2=1.72
r41 9 15 2.79298 $w=4.23e-07 $l=1.03e-07 $layer=LI1_cond $X=6.902 $Y=1.932
+ $X2=6.902 $Y2=2.035
r42 9 11 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=6.902 $Y=1.932
+ $X2=6.902 $Y2=1.885
r43 2 26 400 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=6.61
+ $Y=1.71 $X2=6.775 $Y2=2.685
r44 2 11 400 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=6.61
+ $Y=1.71 $X2=6.775 $Y2=1.885
r45 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.595
+ $Y=0.37 $X2=6.735 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%Q_N 1 2 9 13 14 15 16 23 32
r18 21 23 1.65126 $w=3.33e-07 $l=4.8e-08 $layer=LI1_cond $X=8.362 $Y=1.987
+ $X2=8.362 $Y2=2.035
r19 15 16 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=8.362 $Y=2.405
+ $X2=8.362 $Y2=2.775
r20 14 21 0.653624 $w=3.33e-07 $l=1.9e-08 $layer=LI1_cond $X=8.362 $Y=1.968
+ $X2=8.362 $Y2=1.987
r21 14 32 7.88131 $w=3.33e-07 $l=1.48e-07 $layer=LI1_cond $X=8.362 $Y=1.968
+ $X2=8.362 $Y2=1.82
r22 14 15 12.1093 $w=3.33e-07 $l=3.52e-07 $layer=LI1_cond $X=8.362 $Y=2.053
+ $X2=8.362 $Y2=2.405
r23 14 23 0.619223 $w=3.33e-07 $l=1.8e-08 $layer=LI1_cond $X=8.362 $Y=2.053
+ $X2=8.362 $Y2=2.035
r24 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.445 $Y=1.13
+ $X2=8.445 $Y2=1.82
r25 7 13 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=8.387 $Y=0.988
+ $X2=8.387 $Y2=1.13
r26 7 9 19.1265 $w=2.83e-07 $l=4.73e-07 $layer=LI1_cond $X=8.387 $Y=0.988
+ $X2=8.387 $Y2=0.515
r27 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=1.985
r28 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.815
r29 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.2 $Y=0.37
+ $X2=8.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBN_1%VGND 1 2 3 4 5 18 24 28 32 37 38 40 41 42 44
+ 49 70 79 80 83 87 93
r91 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r92 87 90 10.8067 $w=5.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.63
+ $Y2=0.515
r93 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r94 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 80 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r96 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r97 77 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=7.91
+ $Y2=0
r98 77 79 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=8.4
+ $Y2=0
r99 76 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r100 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r101 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r102 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r103 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r104 70 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.91
+ $Y2=0
r105 70 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r106 69 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r107 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r108 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r109 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r110 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r111 63 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r112 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r113 60 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r114 59 62 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r115 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r116 57 87 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.63
+ $Y2=0
r117 57 59 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.915 $Y=0
+ $X2=3.12 $Y2=0
r118 56 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r119 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r120 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r121 53 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r122 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r123 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r124 50 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.795
+ $Y2=0
r125 50 52 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r126 49 87 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.63
+ $Y2=0
r127 49 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.345 $Y=0
+ $X2=2.16 $Y2=0
r128 47 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r129 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r130 44 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.795
+ $Y2=0
r131 44 46 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r132 42 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r133 42 60 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=3.12
+ $Y2=0
r134 40 68 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=6.03 $Y=0 $X2=6 $Y2=0
r135 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.03 $Y=0 $X2=6.195
+ $Y2=0
r136 39 72 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.36 $Y=0 $X2=6.48
+ $Y2=0
r137 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.36 $Y=0 $X2=6.195
+ $Y2=0
r138 37 62 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.56
+ $Y2=0
r139 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.855
+ $Y2=0
r140 36 65 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.98 $Y=0 $X2=5.04
+ $Y2=0
r141 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.98 $Y=0 $X2=4.855
+ $Y2=0
r142 32 34 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=7.91 $Y=0.495
+ $X2=7.91 $Y2=0.965
r143 30 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r144 30 32 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.495
r145 26 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=0.085
+ $X2=6.195 $Y2=0
r146 26 28 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.195 $Y=0.085
+ $X2=6.195 $Y2=0.495
r147 22 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=0.085
+ $X2=4.855 $Y2=0
r148 22 24 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=4.855 $Y=0.085
+ $X2=4.855 $Y2=0.8
r149 18 20 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.795 $Y=0.515
+ $X2=0.795 $Y2=0.925
r150 16 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r151 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.515
r152 5 34 182 $w=1.7e-07 $l=5.05124e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.56 $X2=7.91 $Y2=0.965
r153 5 32 182 $w=1.7e-07 $l=2.55441e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.56 $X2=7.91 $Y2=0.495
r154 4 28 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.055
+ $Y=0.37 $X2=6.195 $Y2=0.495
r155 3 24 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=4.595
+ $Y=0.59 $X2=4.815 $Y2=0.8
r156 2 90 182 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.37 $X2=2.63 $Y2=0.515
r157 1 20 182 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.56 $X2=0.795 $Y2=0.925
r158 1 18 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.56 $X2=0.795 $Y2=0.515
.ends

