* File: sky130_fd_sc_hs__a221o_4.pxi.spice
* Created: Thu Aug 27 20:25:49 2020
* 
x_PM_SKY130_FD_SC_HS__A221O_4%A1 N_A1_M1005_g N_A1_c_160_n N_A1_c_161_n
+ N_A1_c_172_n N_A1_M1001_g N_A1_c_162_n N_A1_c_163_n N_A1_M1007_g N_A1_c_165_n
+ N_A1_c_166_n N_A1_c_167_n N_A1_c_174_n N_A1_M1004_g N_A1_c_168_n A1 A1
+ N_A1_c_170_n PM_SKY130_FD_SC_HS__A221O_4%A1
x_PM_SKY130_FD_SC_HS__A221O_4%A2 N_A2_c_232_n N_A2_c_240_n N_A2_M1013_g
+ N_A2_M1022_g N_A2_c_234_n N_A2_c_242_n N_A2_M1015_g N_A2_c_235_n N_A2_M1027_g
+ N_A2_c_236_n A2 N_A2_c_238_n PM_SKY130_FD_SC_HS__A221O_4%A2
x_PM_SKY130_FD_SC_HS__A221O_4%A_154_135# N_A_154_135#_M1005_d
+ N_A_154_135#_M1024_d N_A_154_135#_M1011_d N_A_154_135#_M1003_d
+ N_A_154_135#_c_317_n N_A_154_135#_M1000_g N_A_154_135#_c_302_n
+ N_A_154_135#_M1002_g N_A_154_135#_c_318_n N_A_154_135#_M1017_g
+ N_A_154_135#_c_303_n N_A_154_135#_M1012_g N_A_154_135#_c_319_n
+ N_A_154_135#_M1019_g N_A_154_135#_c_304_n N_A_154_135#_M1020_g
+ N_A_154_135#_c_320_n N_A_154_135#_M1025_g N_A_154_135#_c_305_n
+ N_A_154_135#_M1023_g N_A_154_135#_c_306_n N_A_154_135#_c_321_n
+ N_A_154_135#_c_307_n N_A_154_135#_c_341_n N_A_154_135#_c_308_n
+ N_A_154_135#_c_309_n N_A_154_135#_c_310_n N_A_154_135#_c_354_p
+ N_A_154_135#_c_311_n N_A_154_135#_c_380_p N_A_154_135#_c_312_n
+ N_A_154_135#_c_313_n N_A_154_135#_c_314_n N_A_154_135#_c_315_n
+ N_A_154_135#_c_316_n PM_SKY130_FD_SC_HS__A221O_4%A_154_135#
x_PM_SKY130_FD_SC_HS__A221O_4%C1 N_C1_M1024_g N_C1_c_517_n N_C1_M1003_g
+ N_C1_M1026_g N_C1_c_514_n N_C1_c_515_n N_C1_c_516_n N_C1_M1006_g C1 C1
+ PM_SKY130_FD_SC_HS__A221O_4%C1
x_PM_SKY130_FD_SC_HS__A221O_4%B2 N_B2_M1014_g N_B2_c_588_n N_B2_M1008_g
+ N_B2_c_577_n N_B2_c_578_n N_B2_M1016_g N_B2_c_590_n N_B2_M1009_g N_B2_c_580_n
+ N_B2_c_581_n N_B2_c_582_n N_B2_c_583_n N_B2_c_584_n N_B2_c_585_n B2
+ N_B2_c_586_n N_B2_c_587_n PM_SKY130_FD_SC_HS__A221O_4%B2
x_PM_SKY130_FD_SC_HS__A221O_4%B1 N_B1_c_678_n N_B1_M1010_g N_B1_M1011_g
+ N_B1_c_679_n N_B1_M1021_g N_B1_M1018_g N_B1_c_675_n B1 B1 N_B1_c_677_n
+ N_B1_c_683_n PM_SKY130_FD_SC_HS__A221O_4%B1
x_PM_SKY130_FD_SC_HS__A221O_4%VPWR N_VPWR_M1001_s N_VPWR_M1004_s N_VPWR_M1015_s
+ N_VPWR_M1017_d N_VPWR_M1025_d N_VPWR_c_724_n N_VPWR_c_725_n N_VPWR_c_726_n
+ N_VPWR_c_727_n N_VPWR_c_728_n N_VPWR_c_729_n N_VPWR_c_730_n N_VPWR_c_731_n
+ N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n VPWR
+ N_VPWR_c_736_n N_VPWR_c_737_n N_VPWR_c_723_n N_VPWR_c_739_n
+ PM_SKY130_FD_SC_HS__A221O_4%VPWR
x_PM_SKY130_FD_SC_HS__A221O_4%A_157_376# N_A_157_376#_M1001_d
+ N_A_157_376#_M1013_d N_A_157_376#_M1008_d N_A_157_376#_M1010_d
+ N_A_157_376#_c_818_n N_A_157_376#_c_812_n N_A_157_376#_c_813_n
+ N_A_157_376#_c_836_n N_A_157_376#_c_814_n N_A_157_376#_c_815_n
+ N_A_157_376#_c_816_n N_A_157_376#_c_856_n N_A_157_376#_c_817_n
+ PM_SKY130_FD_SC_HS__A221O_4%A_157_376#
x_PM_SKY130_FD_SC_HS__A221O_4%X N_X_M1002_d N_X_M1020_d N_X_M1000_s N_X_M1019_s
+ N_X_c_910_n N_X_c_922_n N_X_c_934_n N_X_c_940_n N_X_c_903_n N_X_c_946_n
+ N_X_c_904_n N_X_c_912_n N_X_c_955_n N_X_c_905_n N_X_c_906_n N_X_c_907_n X
+ N_X_c_909_n PM_SKY130_FD_SC_HS__A221O_4%X
x_PM_SKY130_FD_SC_HS__A221O_4%A_1102_392# N_A_1102_392#_M1003_s
+ N_A_1102_392#_M1006_s N_A_1102_392#_M1009_s N_A_1102_392#_M1021_s
+ N_A_1102_392#_c_1024_n N_A_1102_392#_c_1025_n N_A_1102_392#_c_1036_n
+ N_A_1102_392#_c_1026_n N_A_1102_392#_c_1027_n N_A_1102_392#_c_1028_n
+ N_A_1102_392#_c_1029_n PM_SKY130_FD_SC_HS__A221O_4%A_1102_392#
x_PM_SKY130_FD_SC_HS__A221O_4%A_71_135# N_A_71_135#_M1005_s N_A_71_135#_M1007_s
+ N_A_71_135#_M1022_d N_A_71_135#_c_1069_n N_A_71_135#_c_1074_n
+ N_A_71_135#_c_1066_n N_A_71_135#_c_1067_n N_A_71_135#_c_1085_n
+ N_A_71_135#_c_1068_n PM_SKY130_FD_SC_HS__A221O_4%A_71_135#
x_PM_SKY130_FD_SC_HS__A221O_4%VGND N_VGND_M1022_s N_VGND_M1027_s N_VGND_M1012_s
+ N_VGND_M1023_s N_VGND_M1026_s N_VGND_M1016_s N_VGND_c_1119_n N_VGND_c_1120_n
+ N_VGND_c_1121_n N_VGND_c_1122_n N_VGND_c_1123_n N_VGND_c_1124_n
+ N_VGND_c_1125_n N_VGND_c_1126_n N_VGND_c_1127_n N_VGND_c_1128_n
+ N_VGND_c_1129_n N_VGND_c_1130_n N_VGND_c_1131_n N_VGND_c_1132_n
+ N_VGND_c_1182_n VGND N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n
+ N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n N_VGND_c_1139_n
+ N_VGND_c_1140_n PM_SKY130_FD_SC_HS__A221O_4%VGND
x_PM_SKY130_FD_SC_HS__A221O_4%A_1346_123# N_A_1346_123#_M1014_d
+ N_A_1346_123#_M1011_s N_A_1346_123#_M1018_s N_A_1346_123#_c_1278_n
+ N_A_1346_123#_c_1261_n N_A_1346_123#_c_1262_n N_A_1346_123#_c_1263_n
+ N_A_1346_123#_c_1264_n N_A_1346_123#_c_1265_n N_A_1346_123#_c_1266_n
+ PM_SKY130_FD_SC_HS__A221O_4%A_1346_123#
cc_1 VNB N_A1_M1005_g 0.0126596f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.995
cc_2 VNB N_A1_c_160_n 0.00582947f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.48
cc_3 VNB N_A1_c_161_n 0.0105088f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.715
cc_4 VNB N_A1_c_162_n 0.0143467f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=0.49
cc_5 VNB N_A1_c_163_n 0.0150623f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=0.49
cc_6 VNB N_A1_M1007_g 0.0108339f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_7 VNB N_A1_c_165_n 0.0202405f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.54
cc_8 VNB N_A1_c_166_n 0.00763938f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.715
cc_9 VNB N_A1_c_167_n 0.0147864f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=0.49
cc_10 VNB N_A1_c_168_n 0.0067715f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.49
cc_11 VNB A1 0.0189889f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_12 VNB N_A1_c_170_n 0.0454186f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.4
cc_13 VNB N_A2_c_232_n 0.0112412f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.39
cc_14 VNB N_A2_M1022_g 0.0102533f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.38
cc_15 VNB N_A2_c_234_n 0.0104206f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=0.49
cc_16 VNB N_A2_c_235_n 0.014937f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_17 VNB N_A2_c_236_n 0.0414269f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_18 VNB A2 0.00844479f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.49
cc_19 VNB N_A2_c_238_n 0.0443821f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.465
cc_20 VNB N_A_154_135#_c_302_n 0.0179122f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.54
cc_21 VNB N_A_154_135#_c_303_n 0.0160784f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_22 VNB N_A_154_135#_c_304_n 0.0162363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_154_135#_c_305_n 0.0189669f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.4
cc_24 VNB N_A_154_135#_c_306_n 3.931e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_154_135#_c_307_n 3.95392e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_154_135#_c_308_n 0.0194191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_154_135#_c_309_n 0.00345068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_154_135#_c_310_n 0.00212477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_154_135#_c_311_n 0.0123759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_154_135#_c_312_n 0.0118988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_154_135#_c_313_n 0.00492041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_154_135#_c_314_n 0.0061434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_154_135#_c_315_n 0.00193979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_154_135#_c_316_n 0.0766303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C1_M1024_g 0.0238103f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.995
cc_36 VNB N_C1_M1026_g 0.0228799f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=0.49
cc_37 VNB N_C1_c_514_n 0.00943777f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.565
cc_38 VNB N_C1_c_515_n 0.0277882f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.39
cc_39 VNB N_C1_c_516_n 0.0157501f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_40 VNB N_B2_c_577_n 0.059418f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.805
cc_41 VNB N_B2_c_578_n 0.0051119f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.38
cc_42 VNB N_B2_M1016_g 0.0282044f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.39
cc_43 VNB N_B2_c_580_n 0.00756482f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.49
cc_44 VNB N_B2_c_581_n 0.0604594f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_45 VNB N_B2_c_582_n 0.00523619f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_46 VNB N_B2_c_583_n 0.00422711f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.465
cc_47 VNB N_B2_c_584_n 0.0139812f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_48 VNB N_B2_c_585_n 0.00620432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_B2_c_586_n 0.0468869f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.49
cc_50 VNB N_B2_c_587_n 0.0168974f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.602
cc_51 VNB N_B1_M1011_g 0.0277209f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.715
cc_52 VNB N_B1_M1018_g 0.0306491f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.39
cc_53 VNB N_B1_c_675_n 0.0346654f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_54 VNB B1 0.035572f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_55 VNB N_B1_c_677_n 0.062292f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.465
cc_56 VNB N_VPWR_c_723_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_X_c_903_n 0.00279061f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.465
cc_58 VNB N_X_c_904_n 0.00252589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_X_c_905_n 0.0161413f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.4
cc_60 VNB N_X_c_906_n 0.0195019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_X_c_907_n 0.0221701f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.565
cc_62 VNB X 0.00470385f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.925
cc_63 VNB N_X_c_909_n 0.00409571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_71_135#_c_1066_n 0.0132978f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.54
cc_65 VNB N_A_71_135#_c_1067_n 8.4331e-19 $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.715
cc_66 VNB N_A_71_135#_c_1068_n 0.0171478f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.49
cc_67 VNB N_VGND_c_1119_n 0.0138474f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.805
cc_68 VNB N_VGND_c_1120_n 0.0162981f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.39
cc_69 VNB N_VGND_c_1121_n 0.0140948f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.465
cc_70 VNB N_VGND_c_1122_n 0.0259638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1123_n 0.0184531f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.4
cc_72 VNB N_VGND_c_1124_n 0.00304657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1125_n 0.0106636f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.602
cc_74 VNB N_VGND_c_1126_n 0.0562111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1127_n 0.00326288f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.41
cc_76 VNB N_VGND_c_1128_n 0.00840773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1129_n 0.0197463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1130_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1131_n 0.0202649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1132_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1133_n 0.022977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1134_n 0.0178473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1135_n 0.0218123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1136_n 0.0572372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1137_n 0.55948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1138_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1139_n 0.013849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1140_n 0.00351416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1346_123#_c_1261_n 0.0126797f $X=-0.19 $Y=-0.245 $X2=1.125
+ $Y2=0.995
cc_90 VNB N_A_1346_123#_c_1262_n 0.00246562f $X=-0.19 $Y=-0.245 $X2=1.125
+ $Y2=0.995
cc_91 VNB N_A_1346_123#_c_1263_n 0.00912157f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.49
cc_92 VNB N_A_1346_123#_c_1264_n 0.0127125f $X=-0.19 $Y=-0.245 $X2=1.28
+ $Y2=1.805
cc_93 VNB N_A_1346_123#_c_1265_n 0.00355281f $X=-0.19 $Y=-0.245 $X2=1.28
+ $Y2=2.38
cc_94 VNB N_A_1346_123#_c_1266_n 0.0255734f $X=-0.19 $Y=-0.245 $X2=1.125
+ $Y2=0.49
cc_95 VPB N_A1_c_161_n 0.00326976f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.715
cc_96 VPB N_A1_c_172_n 0.0238538f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.805
cc_97 VPB N_A1_c_166_n 0.00325983f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=1.715
cc_98 VPB N_A1_c_174_n 0.0249695f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=1.805
cc_99 VPB N_A2_c_232_n 0.00302156f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.39
cc_100 VPB N_A2_c_240_n 0.0236606f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=0.995
cc_101 VPB N_A2_c_234_n 0.00275598f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=0.49
cc_102 VPB N_A2_c_242_n 0.0219214f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.565
cc_103 VPB N_A_154_135#_c_317_n 0.0170281f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.39
cc_104 VPB N_A_154_135#_c_318_n 0.0151113f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0.49
cc_105 VPB N_A_154_135#_c_319_n 0.0151113f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.465
cc_106 VPB N_A_154_135#_c_320_n 0.0191176f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_154_135#_c_321_n 0.00260596f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0.925
cc_108 VPB N_A_154_135#_c_307_n 0.00563034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_154_135#_c_311_n 0.0099801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_154_135#_c_312_n 0.0181036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_154_135#_c_313_n 0.00399505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_154_135#_c_316_n 0.0482838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_C1_c_517_n 0.0167242f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.48
cc_114 VPB N_C1_c_515_n 0.0314573f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.39
cc_115 VPB N_C1_c_516_n 0.0262421f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.995
cc_116 VPB C1 0.0157039f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=0.49
cc_117 VPB N_B2_c_588_n 0.0148151f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=0.995
cc_118 VPB N_B2_c_578_n 0.00543929f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=2.38
cc_119 VPB N_B2_c_590_n 0.0163552f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.995
cc_120 VPB N_B2_c_582_n 0.0105237f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.38
cc_121 VPB N_B2_c_583_n 0.0253291f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.465
cc_122 VPB N_B1_c_678_n 0.0166636f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=0.565
cc_123 VPB N_B1_c_679_n 0.0186548f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=2.38
cc_124 VPB N_B1_c_675_n 0.0415078f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.995
cc_125 VPB B1 0.019573f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.38
cc_126 VPB N_B1_c_677_n 0.026591f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.465
cc_127 VPB N_B1_c_683_n 0.0125041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_724_n 0.0410772f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=0.49
cc_129 VPB N_VPWR_c_725_n 0.00894283f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.38
cc_130 VPB N_VPWR_c_726_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_727_n 0.0113661f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=0.84
cc_132 VPB N_VPWR_c_728_n 0.0123263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_729_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.4
cc_134 VPB N_VPWR_c_730_n 0.0225995f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.4
cc_135 VPB N_VPWR_c_731_n 0.00614296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_732_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_733_n 0.00601813f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0.565
cc_138 VPB N_VPWR_c_734_n 0.0177589f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0.925
cc_139 VPB N_VPWR_c_735_n 0.00613001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_736_n 0.0214857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_737_n 0.116915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_723_n 0.138173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_739_n 0.0346291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_157_376#_c_812_n 0.0295027f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0.49
cc_145 VPB N_A_157_376#_c_813_n 0.00183108f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.38
cc_146 VPB N_A_157_376#_c_814_n 0.00439731f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.39
cc_147 VPB N_A_157_376#_c_815_n 0.00330685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_157_376#_c_816_n 0.00293822f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=0.84
cc_149 VPB N_A_157_376#_c_817_n 0.00212467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_X_c_910_n 0.016621f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.995
cc_151 VPB N_X_c_907_n 0.0140119f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0.565
cc_152 VPB N_A_1102_392#_c_1024_n 0.0122177f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.39
cc_153 VPB N_A_1102_392#_c_1025_n 0.00312572f $X=-0.19 $Y=1.66 $X2=1.28
+ $Y2=1.715
cc_154 VPB N_A_1102_392#_c_1026_n 0.013123f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.39
cc_155 VPB N_A_1102_392#_c_1027_n 0.0381703f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=1.465
cc_156 VPB N_A_1102_392#_c_1028_n 0.00124149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_1102_392#_c_1029_n 0.00338059f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.4
cc_158 N_A1_c_166_n N_A2_c_232_n 0.00232278f $X=1.28 $Y=1.715 $X2=0 $Y2=0
cc_159 N_A1_c_174_n N_A2_c_240_n 0.00232278f $X=1.28 $Y=1.805 $X2=0 $Y2=0
cc_160 N_A1_c_170_n N_A2_M1022_g 7.29007e-19 $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_161 N_A1_c_165_n N_A2_c_236_n 0.00232278f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_162 N_A1_c_170_n N_A2_c_238_n 0.00509489f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_163 N_A1_M1005_g N_A_154_135#_c_306_n 0.00834817f $X=0.695 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A1_c_160_n N_A_154_135#_c_306_n 0.0033001f $X=0.71 $Y=1.48 $X2=0 $Y2=0
cc_165 N_A1_c_161_n N_A_154_135#_c_306_n 0.00299664f $X=0.71 $Y=1.715 $X2=0
+ $Y2=0
cc_166 N_A1_M1007_g N_A_154_135#_c_306_n 0.00409333f $X=1.125 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A1_c_165_n N_A_154_135#_c_306_n 0.00830365f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_168 N_A1_c_166_n N_A_154_135#_c_306_n 0.0010381f $X=1.28 $Y=1.715 $X2=0 $Y2=0
cc_169 N_A1_c_161_n N_A_154_135#_c_321_n 0.00464588f $X=0.71 $Y=1.715 $X2=0
+ $Y2=0
cc_170 N_A1_c_172_n N_A_154_135#_c_321_n 0.0018759f $X=0.71 $Y=1.805 $X2=0 $Y2=0
cc_171 N_A1_c_165_n N_A_154_135#_c_312_n 0.0042433f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_172 N_A1_c_166_n N_A_154_135#_c_312_n 0.00992585f $X=1.28 $Y=1.715 $X2=0
+ $Y2=0
cc_173 N_A1_c_174_n N_A_154_135#_c_312_n 0.00406102f $X=1.28 $Y=1.805 $X2=0
+ $Y2=0
cc_174 N_A1_c_172_n N_VPWR_c_724_n 0.0125171f $X=0.71 $Y=1.805 $X2=0 $Y2=0
cc_175 N_A1_c_174_n N_VPWR_c_724_n 6.83173e-19 $X=1.28 $Y=1.805 $X2=0 $Y2=0
cc_176 N_A1_c_172_n N_VPWR_c_736_n 0.00467292f $X=0.71 $Y=1.805 $X2=0 $Y2=0
cc_177 N_A1_c_174_n N_VPWR_c_736_n 0.00507376f $X=1.28 $Y=1.805 $X2=0 $Y2=0
cc_178 N_A1_c_172_n N_VPWR_c_723_n 0.00471987f $X=0.71 $Y=1.805 $X2=0 $Y2=0
cc_179 N_A1_c_174_n N_VPWR_c_723_n 0.00520574f $X=1.28 $Y=1.805 $X2=0 $Y2=0
cc_180 N_A1_c_174_n N_VPWR_c_739_n 0.011073f $X=1.28 $Y=1.805 $X2=0 $Y2=0
cc_181 N_A1_c_174_n N_A_157_376#_c_818_n 0.0136739f $X=1.28 $Y=1.805 $X2=0 $Y2=0
cc_182 N_A1_c_172_n N_A_157_376#_c_815_n 0.00613047f $X=0.71 $Y=1.805 $X2=0
+ $Y2=0
cc_183 N_A1_c_174_n N_A_157_376#_c_815_n 0.0113213f $X=1.28 $Y=1.805 $X2=0 $Y2=0
cc_184 N_A1_c_172_n N_X_c_912_n 0.0181906f $X=0.71 $Y=1.805 $X2=0 $Y2=0
cc_185 N_A1_c_165_n N_X_c_912_n 2.3069e-19 $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_186 N_A1_c_174_n N_X_c_912_n 0.0132438f $X=1.28 $Y=1.805 $X2=0 $Y2=0
cc_187 N_A1_M1005_g N_X_c_905_n 0.00523379f $X=0.695 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_M1007_g N_X_c_905_n 0.00454499f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_165_n N_X_c_905_n 0.00165477f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_190 A1 N_X_c_905_n 0.00437127f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_191 N_A1_M1005_g N_X_c_906_n 0.00206546f $X=0.695 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_M1005_g N_X_c_907_n 0.0122199f $X=0.695 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A1_c_172_n N_X_c_907_n 0.00359625f $X=0.71 $Y=1.805 $X2=0 $Y2=0
cc_194 N_A1_M1005_g N_A_71_135#_c_1069_n 0.0102992f $X=0.695 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A1_c_162_n N_A_71_135#_c_1069_n 0.00238533f $X=1.05 $Y=0.49 $X2=0 $Y2=0
cc_196 N_A1_M1007_g N_A_71_135#_c_1069_n 0.0131077f $X=1.125 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A1_c_167_n N_A_71_135#_c_1069_n 0.00448161f $X=1.435 $Y=0.49 $X2=0
+ $Y2=0
cc_198 A1 N_A_71_135#_c_1069_n 0.0140569f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_199 A1 N_A_71_135#_c_1074_n 0.00994896f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_200 N_A1_c_167_n N_A_71_135#_c_1066_n 0.00234729f $X=1.435 $Y=0.49 $X2=0
+ $Y2=0
cc_201 A1 N_A_71_135#_c_1066_n 0.0131478f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_202 N_A1_c_170_n N_A_71_135#_c_1066_n 3.82631e-19 $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_203 N_A1_M1007_g N_A_71_135#_c_1067_n 0.00288366f $X=1.125 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A1_c_165_n N_A_71_135#_c_1067_n 0.00529894f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_205 N_A1_M1005_g N_A_71_135#_c_1068_n 7.91278e-19 $X=0.695 $Y=0.995 $X2=0
+ $Y2=0
cc_206 A1 N_VGND_c_1119_n 0.0315455f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_207 N_A1_c_170_n N_VGND_c_1119_n 0.00162808f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_208 N_A1_c_163_n N_VGND_c_1126_n 0.0175556f $X=0.77 $Y=0.49 $X2=0 $Y2=0
cc_209 A1 N_VGND_c_1126_n 0.021134f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_210 N_A1_c_170_n N_VGND_c_1126_n 0.0056689f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_211 A1 N_VGND_c_1128_n 0.0294117f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_212 N_A1_c_163_n N_VGND_c_1137_n 0.0244466f $X=0.77 $Y=0.49 $X2=0 $Y2=0
cc_213 A1 N_VGND_c_1137_n 0.011067f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_214 N_A1_c_170_n N_VGND_c_1137_n 0.00759015f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_215 N_A2_c_242_n N_A_154_135#_c_317_n 0.0266739f $X=2.625 $Y=1.805 $X2=0
+ $Y2=0
cc_216 N_A2_c_235_n N_A_154_135#_c_302_n 0.0131106f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_217 N_A2_c_238_n N_A_154_135#_c_302_n 0.00102307f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_218 N_A2_c_236_n N_A_154_135#_c_341_n 3.22675e-19 $X=2.89 $Y=1.405 $X2=0
+ $Y2=0
cc_219 N_A2_c_232_n N_A_154_135#_c_312_n 0.00895806f $X=2.175 $Y=1.715 $X2=0
+ $Y2=0
cc_220 N_A2_c_240_n N_A_154_135#_c_312_n 0.0039296f $X=2.175 $Y=1.805 $X2=0
+ $Y2=0
cc_221 N_A2_c_234_n N_A_154_135#_c_312_n 0.00839595f $X=2.625 $Y=1.715 $X2=0
+ $Y2=0
cc_222 N_A2_c_242_n N_A_154_135#_c_312_n 0.00377824f $X=2.625 $Y=1.805 $X2=0
+ $Y2=0
cc_223 N_A2_c_236_n N_A_154_135#_c_312_n 0.0127287f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_224 N_A2_c_234_n N_A_154_135#_c_316_n 0.00733989f $X=2.625 $Y=1.715 $X2=0
+ $Y2=0
cc_225 N_A2_c_236_n N_A_154_135#_c_316_n 0.0131106f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_226 N_A2_c_242_n N_VPWR_c_725_n 0.00479437f $X=2.625 $Y=1.805 $X2=0 $Y2=0
cc_227 N_A2_c_240_n N_VPWR_c_730_n 0.00507376f $X=2.175 $Y=1.805 $X2=0 $Y2=0
cc_228 N_A2_c_242_n N_VPWR_c_730_n 0.00507376f $X=2.625 $Y=1.805 $X2=0 $Y2=0
cc_229 N_A2_c_240_n N_VPWR_c_723_n 0.00520574f $X=2.175 $Y=1.805 $X2=0 $Y2=0
cc_230 N_A2_c_242_n N_VPWR_c_723_n 0.00520574f $X=2.625 $Y=1.805 $X2=0 $Y2=0
cc_231 N_A2_c_240_n N_VPWR_c_739_n 0.0111326f $X=2.175 $Y=1.805 $X2=0 $Y2=0
cc_232 N_A2_c_240_n N_A_157_376#_c_818_n 0.0136739f $X=2.175 $Y=1.805 $X2=0
+ $Y2=0
cc_233 N_A2_c_242_n N_A_157_376#_c_812_n 0.0102143f $X=2.625 $Y=1.805 $X2=0
+ $Y2=0
cc_234 N_A2_c_240_n N_A_157_376#_c_816_n 0.0116249f $X=2.175 $Y=1.805 $X2=0
+ $Y2=0
cc_235 N_A2_c_242_n N_A_157_376#_c_816_n 0.00915684f $X=2.625 $Y=1.805 $X2=0
+ $Y2=0
cc_236 N_A2_c_242_n N_X_c_922_n 0.00297598f $X=2.625 $Y=1.805 $X2=0 $Y2=0
cc_237 N_A2_c_235_n N_X_c_903_n 6.23275e-19 $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_238 N_A2_c_240_n N_X_c_912_n 0.0126447f $X=2.175 $Y=1.805 $X2=0 $Y2=0
cc_239 N_A2_c_242_n N_X_c_912_n 0.0119302f $X=2.625 $Y=1.805 $X2=0 $Y2=0
cc_240 N_A2_M1022_g N_X_c_905_n 0.00540271f $X=2.46 $Y=0.935 $X2=0 $Y2=0
cc_241 N_A2_c_235_n N_X_c_905_n 0.00725658f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_242 N_A2_c_236_n N_X_c_905_n 0.00189607f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_243 A2 N_X_c_905_n 8.85114e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_244 N_A2_c_235_n X 7.93272e-19 $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_245 N_A2_c_236_n X 8.83029e-19 $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_246 N_A2_c_235_n N_X_c_909_n 0.00276942f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_247 A2 N_A_71_135#_M1022_d 0.00219033f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_248 N_A2_M1022_g N_A_71_135#_c_1066_n 0.0070549f $X=2.46 $Y=0.935 $X2=0 $Y2=0
cc_249 N_A2_c_235_n N_A_71_135#_c_1066_n 6.08595e-19 $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_250 N_A2_c_236_n N_A_71_135#_c_1066_n 0.0231609f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_251 N_A2_M1022_g N_A_71_135#_c_1085_n 0.00996461f $X=2.46 $Y=0.935 $X2=0
+ $Y2=0
cc_252 A2 N_A_71_135#_c_1085_n 0.0145781f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_253 N_A2_c_238_n N_A_71_135#_c_1085_n 2.47224e-19 $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_254 N_A2_M1022_g N_VGND_c_1119_n 0.00270215f $X=2.46 $Y=0.935 $X2=0 $Y2=0
cc_255 A2 N_VGND_c_1119_n 0.0255727f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_256 N_A2_c_238_n N_VGND_c_1119_n 0.00308142f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_257 N_A2_c_235_n N_VGND_c_1120_n 0.00240899f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_258 A2 N_VGND_c_1120_n 0.0246703f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_259 N_A2_c_238_n N_VGND_c_1120_n 0.00262568f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_260 N_A2_c_236_n N_VGND_c_1128_n 0.00144271f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_261 A2 N_VGND_c_1128_n 0.0039865f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_262 N_A2_c_238_n N_VGND_c_1128_n 4.08097e-19 $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_263 N_A2_c_235_n N_VGND_c_1133_n 0.00420632f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_264 A2 N_VGND_c_1133_n 0.0315176f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_265 N_A2_c_238_n N_VGND_c_1133_n 0.00659434f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_266 N_A2_c_235_n N_VGND_c_1137_n 0.00472204f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_267 A2 N_VGND_c_1137_n 0.0168113f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_268 N_A2_c_238_n N_VGND_c_1137_n 0.0103546f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_269 N_A_154_135#_c_308_n N_C1_M1024_g 0.0128795f $X=5.61 $Y=1.215 $X2=0 $Y2=0
cc_270 N_A_154_135#_c_309_n N_C1_M1024_g 0.0119691f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_271 N_A_154_135#_c_310_n N_C1_M1024_g 8.66403e-19 $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_272 N_A_154_135#_c_313_n N_C1_M1024_g 0.00339201f $X=4.795 $Y=1.215 $X2=0
+ $Y2=0
cc_273 N_A_154_135#_c_314_n N_C1_M1024_g 0.00142589f $X=5.85 $Y=1.215 $X2=0
+ $Y2=0
cc_274 N_A_154_135#_c_354_p N_C1_c_517_n 0.00555346f $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_275 N_A_154_135#_c_309_n N_C1_M1026_g 0.00714623f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_276 N_A_154_135#_c_310_n N_C1_M1026_g 0.00509715f $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_277 N_A_154_135#_c_314_n N_C1_M1026_g 0.0109783f $X=5.85 $Y=1.215 $X2=0 $Y2=0
cc_278 N_A_154_135#_c_310_n N_C1_c_514_n 0.00730338f $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_279 N_A_154_135#_c_315_n N_C1_c_514_n 0.00190788f $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_280 N_A_154_135#_c_308_n N_C1_c_515_n 0.00190609f $X=5.61 $Y=1.215 $X2=0
+ $Y2=0
cc_281 N_A_154_135#_c_310_n N_C1_c_515_n 0.00580359f $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_282 N_A_154_135#_c_354_p N_C1_c_515_n 0.00316755f $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_283 N_A_154_135#_c_313_n N_C1_c_515_n 0.00556938f $X=4.795 $Y=1.215 $X2=0
+ $Y2=0
cc_284 N_A_154_135#_c_314_n N_C1_c_515_n 0.00459898f $X=5.85 $Y=1.215 $X2=0
+ $Y2=0
cc_285 N_A_154_135#_c_315_n N_C1_c_515_n 0.00502274f $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_286 N_A_154_135#_c_316_n N_C1_c_515_n 8.07662e-19 $X=4.585 $Y=1.557 $X2=0
+ $Y2=0
cc_287 N_A_154_135#_c_354_p N_C1_c_516_n 0.0102662f $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_288 N_A_154_135#_c_311_n N_C1_c_516_n 0.0104813f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_289 N_A_154_135#_c_315_n N_C1_c_516_n 0.00303754f $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_290 N_A_154_135#_c_308_n C1 0.015801f $X=5.61 $Y=1.215 $X2=0 $Y2=0
cc_291 N_A_154_135#_c_310_n C1 0.00864364f $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_292 N_A_154_135#_c_354_p C1 0.0205379f $X=6.085 $Y=2.105 $X2=0 $Y2=0
cc_293 N_A_154_135#_c_313_n C1 0.00900014f $X=4.795 $Y=1.215 $X2=0 $Y2=0
cc_294 N_A_154_135#_c_314_n C1 0.0109932f $X=5.85 $Y=1.215 $X2=0 $Y2=0
cc_295 N_A_154_135#_c_315_n C1 0.0126759f $X=6.085 $Y=1.685 $X2=0 $Y2=0
cc_296 N_A_154_135#_c_354_p N_B2_c_588_n 9.94577e-19 $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_297 N_A_154_135#_c_311_n N_B2_c_578_n 0.00518731f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_298 N_A_154_135#_c_311_n N_B2_M1016_g 0.00307374f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_299 N_A_154_135#_c_311_n N_B2_c_580_n 0.00290892f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_300 N_A_154_135#_c_380_p N_B2_c_580_n 5.1726e-19 $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_301 N_A_154_135#_c_380_p N_B2_c_581_n 2.91453e-19 $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_302 N_A_154_135#_c_354_p N_B2_c_582_n 5.48709e-19 $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_303 N_A_154_135#_c_311_n N_B2_c_582_n 0.0102511f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_304 N_A_154_135#_c_311_n N_B2_c_583_n 0.0141302f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_305 N_A_154_135#_c_311_n N_B2_c_584_n 0.00279407f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_306 N_A_154_135#_c_380_p N_B2_c_584_n 2.5461e-19 $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_307 N_A_154_135#_c_310_n N_B2_c_587_n 5.938e-19 $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_308 N_A_154_135#_c_311_n N_B2_c_587_n 0.00433746f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_309 N_A_154_135#_c_314_n N_B2_c_587_n 2.42029e-19 $X=5.85 $Y=1.215 $X2=0
+ $Y2=0
cc_310 N_A_154_135#_c_380_p N_B1_M1011_g 0.0136043f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_311 N_A_154_135#_c_380_p N_B1_M1018_g 0.0186666f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_312 N_A_154_135#_c_311_n N_B1_c_675_n 0.032731f $X=8.115 $Y=1.685 $X2=0 $Y2=0
cc_313 N_A_154_135#_c_380_p N_B1_c_675_n 0.0180239f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_314 N_A_154_135#_c_380_p B1 0.00257795f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_315 N_A_154_135#_c_311_n N_B1_c_683_n 0.0127433f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_316 N_A_154_135#_c_380_p N_B1_c_683_n 0.0238299f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_317 N_A_154_135#_c_317_n N_VPWR_c_725_n 0.0096174f $X=3.235 $Y=1.765 $X2=0
+ $Y2=0
cc_318 N_A_154_135#_c_318_n N_VPWR_c_725_n 0.00115327f $X=3.685 $Y=1.765 $X2=0
+ $Y2=0
cc_319 N_A_154_135#_c_317_n N_VPWR_c_726_n 0.00115327f $X=3.235 $Y=1.765 $X2=0
+ $Y2=0
cc_320 N_A_154_135#_c_318_n N_VPWR_c_726_n 0.0089303f $X=3.685 $Y=1.765 $X2=0
+ $Y2=0
cc_321 N_A_154_135#_c_319_n N_VPWR_c_726_n 0.0089303f $X=4.135 $Y=1.765 $X2=0
+ $Y2=0
cc_322 N_A_154_135#_c_320_n N_VPWR_c_726_n 0.00115327f $X=4.585 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A_154_135#_c_319_n N_VPWR_c_727_n 0.00115327f $X=4.135 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_A_154_135#_c_320_n N_VPWR_c_727_n 0.00992118f $X=4.585 $Y=1.765 $X2=0
+ $Y2=0
cc_325 N_A_154_135#_c_317_n N_VPWR_c_732_n 0.00413917f $X=3.235 $Y=1.765 $X2=0
+ $Y2=0
cc_326 N_A_154_135#_c_318_n N_VPWR_c_732_n 0.00413917f $X=3.685 $Y=1.765 $X2=0
+ $Y2=0
cc_327 N_A_154_135#_c_319_n N_VPWR_c_734_n 0.00413917f $X=4.135 $Y=1.765 $X2=0
+ $Y2=0
cc_328 N_A_154_135#_c_320_n N_VPWR_c_734_n 0.00413917f $X=4.585 $Y=1.765 $X2=0
+ $Y2=0
cc_329 N_A_154_135#_c_317_n N_VPWR_c_723_n 0.00405449f $X=3.235 $Y=1.765 $X2=0
+ $Y2=0
cc_330 N_A_154_135#_c_318_n N_VPWR_c_723_n 0.00405449f $X=3.685 $Y=1.765 $X2=0
+ $Y2=0
cc_331 N_A_154_135#_c_319_n N_VPWR_c_723_n 0.00405449f $X=4.135 $Y=1.765 $X2=0
+ $Y2=0
cc_332 N_A_154_135#_c_320_n N_VPWR_c_723_n 0.00405449f $X=4.585 $Y=1.765 $X2=0
+ $Y2=0
cc_333 N_A_154_135#_M1003_d N_A_157_376#_c_812_n 0.0039258f $X=5.935 $Y=1.96
+ $X2=0 $Y2=0
cc_334 N_A_154_135#_c_317_n N_A_157_376#_c_812_n 0.0125709f $X=3.235 $Y=1.765
+ $X2=0 $Y2=0
cc_335 N_A_154_135#_c_318_n N_A_157_376#_c_812_n 0.0118864f $X=3.685 $Y=1.765
+ $X2=0 $Y2=0
cc_336 N_A_154_135#_c_319_n N_A_157_376#_c_812_n 0.0118864f $X=4.135 $Y=1.765
+ $X2=0 $Y2=0
cc_337 N_A_154_135#_c_320_n N_A_157_376#_c_812_n 0.0156754f $X=4.585 $Y=1.765
+ $X2=0 $Y2=0
cc_338 N_A_154_135#_c_307_n N_A_157_376#_c_812_n 0.00421634f $X=4.71 $Y=1.55
+ $X2=0 $Y2=0
cc_339 N_A_154_135#_c_354_p N_A_157_376#_c_812_n 0.0170874f $X=6.085 $Y=2.105
+ $X2=0 $Y2=0
cc_340 N_A_154_135#_c_311_n N_A_157_376#_c_812_n 0.0138383f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_341 N_A_154_135#_c_313_n N_A_157_376#_c_812_n 0.00543313f $X=4.795 $Y=1.215
+ $X2=0 $Y2=0
cc_342 N_A_154_135#_c_354_p N_A_157_376#_c_813_n 0.00499324f $X=6.085 $Y=2.105
+ $X2=0 $Y2=0
cc_343 N_A_154_135#_c_311_n N_A_157_376#_c_813_n 0.0263738f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_344 N_A_154_135#_c_354_p N_A_157_376#_c_836_n 0.00220216f $X=6.085 $Y=2.105
+ $X2=0 $Y2=0
cc_345 N_A_154_135#_c_311_n N_A_157_376#_c_814_n 0.0616025f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_346 N_A_154_135#_c_317_n N_A_157_376#_c_816_n 9.48742e-19 $X=3.235 $Y=1.765
+ $X2=0 $Y2=0
cc_347 N_A_154_135#_c_311_n N_A_157_376#_c_817_n 0.0332709f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_348 N_A_154_135#_c_341_n N_X_c_922_n 0.0752512f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_349 N_A_154_135#_c_317_n N_X_c_934_n 0.0120803f $X=3.235 $Y=1.765 $X2=0 $Y2=0
cc_350 N_A_154_135#_c_318_n N_X_c_934_n 0.0113147f $X=3.685 $Y=1.765 $X2=0 $Y2=0
cc_351 N_A_154_135#_c_319_n N_X_c_934_n 0.0113147f $X=4.135 $Y=1.765 $X2=0 $Y2=0
cc_352 N_A_154_135#_c_320_n N_X_c_934_n 0.0127916f $X=4.585 $Y=1.765 $X2=0 $Y2=0
cc_353 N_A_154_135#_c_307_n N_X_c_934_n 0.0752512f $X=4.71 $Y=1.55 $X2=0 $Y2=0
cc_354 N_A_154_135#_c_316_n N_X_c_934_n 0.00447689f $X=4.585 $Y=1.557 $X2=0
+ $Y2=0
cc_355 N_A_154_135#_c_302_n N_X_c_940_n 0.0110688f $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_356 N_A_154_135#_c_312_n N_X_c_940_n 0.00529375f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_357 N_A_154_135#_c_316_n N_X_c_940_n 0.0014255f $X=4.585 $Y=1.557 $X2=0 $Y2=0
cc_358 N_A_154_135#_c_302_n N_X_c_903_n 0.0085362f $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_359 N_A_154_135#_c_303_n N_X_c_903_n 0.00805676f $X=3.81 $Y=1.35 $X2=0 $Y2=0
cc_360 N_A_154_135#_c_304_n N_X_c_903_n 5.86626e-19 $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_361 N_A_154_135#_c_303_n N_X_c_946_n 0.0109154f $X=3.81 $Y=1.35 $X2=0 $Y2=0
cc_362 N_A_154_135#_c_304_n N_X_c_946_n 0.01168f $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_363 N_A_154_135#_c_307_n N_X_c_946_n 0.0182043f $X=4.71 $Y=1.55 $X2=0 $Y2=0
cc_364 N_A_154_135#_c_341_n N_X_c_946_n 0.0348755f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_365 N_A_154_135#_c_316_n N_X_c_946_n 0.00467805f $X=4.585 $Y=1.557 $X2=0
+ $Y2=0
cc_366 N_A_154_135#_c_303_n N_X_c_904_n 5.76374e-19 $X=3.81 $Y=1.35 $X2=0 $Y2=0
cc_367 N_A_154_135#_c_304_n N_X_c_904_n 0.00715462f $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_368 N_A_154_135#_c_321_n N_X_c_912_n 0.0244299f $X=1.075 $Y=1.665 $X2=0 $Y2=0
cc_369 N_A_154_135#_c_312_n N_X_c_912_n 0.0752512f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_370 N_A_154_135#_c_302_n N_X_c_955_n 9.42568e-19 $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_371 N_A_154_135#_c_303_n N_X_c_955_n 7.32094e-19 $X=3.81 $Y=1.35 $X2=0 $Y2=0
cc_372 N_A_154_135#_c_341_n N_X_c_955_n 0.0111425f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_373 N_A_154_135#_c_312_n N_X_c_955_n 0.00527902f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_374 N_A_154_135#_c_316_n N_X_c_955_n 0.00266594f $X=4.585 $Y=1.557 $X2=0
+ $Y2=0
cc_375 N_A_154_135#_c_306_n N_X_c_905_n 0.0195291f $X=0.91 $Y=1.165 $X2=0 $Y2=0
cc_376 N_A_154_135#_c_312_n N_X_c_905_n 0.0235768f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_377 N_A_154_135#_c_306_n N_X_c_906_n 0.0022879f $X=0.91 $Y=1.165 $X2=0 $Y2=0
cc_378 N_A_154_135#_c_306_n N_X_c_907_n 0.0132312f $X=0.91 $Y=1.165 $X2=0 $Y2=0
cc_379 N_A_154_135#_c_321_n N_X_c_907_n 0.00741348f $X=1.075 $Y=1.665 $X2=0
+ $Y2=0
cc_380 N_A_154_135#_c_302_n X 0.0047024f $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_381 N_A_154_135#_c_341_n X 0.00163342f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_382 N_A_154_135#_c_312_n X 0.00413468f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_383 N_A_154_135#_c_316_n X 9.39344e-19 $X=4.585 $Y=1.557 $X2=0 $Y2=0
cc_384 N_A_154_135#_c_302_n N_X_c_909_n 0.00476106f $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_385 N_A_154_135#_c_341_n N_X_c_909_n 0.00184559f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_386 N_A_154_135#_c_312_n N_X_c_909_n 0.015136f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_387 N_A_154_135#_c_316_n N_X_c_909_n 0.00169047f $X=4.585 $Y=1.557 $X2=0
+ $Y2=0
cc_388 N_A_154_135#_M1003_d N_A_1102_392#_c_1024_n 0.00203088f $X=5.935 $Y=1.96
+ $X2=0 $Y2=0
cc_389 N_A_154_135#_M1005_d N_A_71_135#_c_1069_n 0.00430941f $X=0.77 $Y=0.675
+ $X2=0 $Y2=0
cc_390 N_A_154_135#_c_306_n N_A_71_135#_c_1069_n 0.0160844f $X=0.91 $Y=1.165
+ $X2=0 $Y2=0
cc_391 N_A_154_135#_c_312_n N_A_71_135#_c_1069_n 0.00136585f $X=3.595 $Y=1.55
+ $X2=0 $Y2=0
cc_392 N_A_154_135#_c_306_n N_A_71_135#_c_1074_n 0.00606866f $X=0.91 $Y=1.165
+ $X2=0 $Y2=0
cc_393 N_A_154_135#_c_312_n N_A_71_135#_c_1066_n 0.0899913f $X=3.595 $Y=1.55
+ $X2=0 $Y2=0
cc_394 N_A_154_135#_c_306_n N_A_71_135#_c_1067_n 0.0104031f $X=0.91 $Y=1.165
+ $X2=0 $Y2=0
cc_395 N_A_154_135#_c_312_n N_A_71_135#_c_1067_n 0.0123781f $X=3.595 $Y=1.55
+ $X2=0 $Y2=0
cc_396 N_A_154_135#_c_308_n N_VGND_M1023_s 0.00837877f $X=5.61 $Y=1.215 $X2=0
+ $Y2=0
cc_397 N_A_154_135#_c_313_n N_VGND_M1023_s 0.00115102f $X=4.795 $Y=1.215 $X2=0
+ $Y2=0
cc_398 N_A_154_135#_c_302_n N_VGND_c_1120_n 0.00278543f $X=3.38 $Y=1.35 $X2=0
+ $Y2=0
cc_399 N_A_154_135#_c_303_n N_VGND_c_1121_n 0.00209581f $X=3.81 $Y=1.35 $X2=0
+ $Y2=0
cc_400 N_A_154_135#_c_304_n N_VGND_c_1121_n 0.00150779f $X=4.24 $Y=1.35 $X2=0
+ $Y2=0
cc_401 N_A_154_135#_c_304_n N_VGND_c_1122_n 4.82085e-19 $X=4.24 $Y=1.35 $X2=0
+ $Y2=0
cc_402 N_A_154_135#_c_305_n N_VGND_c_1122_n 0.0133684f $X=4.67 $Y=1.35 $X2=0
+ $Y2=0
cc_403 N_A_154_135#_c_308_n N_VGND_c_1122_n 0.0445845f $X=5.61 $Y=1.215 $X2=0
+ $Y2=0
cc_404 N_A_154_135#_c_309_n N_VGND_c_1122_n 0.0151478f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_405 N_A_154_135#_c_313_n N_VGND_c_1122_n 0.00887034f $X=4.795 $Y=1.215 $X2=0
+ $Y2=0
cc_406 N_A_154_135#_c_309_n N_VGND_c_1123_n 0.00646413f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_407 N_A_154_135#_c_309_n N_VGND_c_1124_n 0.00765349f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_408 N_A_154_135#_c_311_n N_VGND_c_1124_n 0.0123214f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_409 N_A_154_135#_c_314_n N_VGND_c_1124_n 0.00721388f $X=5.85 $Y=1.215 $X2=0
+ $Y2=0
cc_410 N_A_154_135#_c_302_n N_VGND_c_1129_n 0.00466874f $X=3.38 $Y=1.35 $X2=0
+ $Y2=0
cc_411 N_A_154_135#_c_303_n N_VGND_c_1129_n 0.00466874f $X=3.81 $Y=1.35 $X2=0
+ $Y2=0
cc_412 N_A_154_135#_c_309_n N_VGND_c_1131_n 0.00739421f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_413 N_A_154_135#_c_309_n N_VGND_c_1182_n 0.020538f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_414 N_A_154_135#_c_311_n N_VGND_c_1182_n 6.72765e-19 $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_415 N_A_154_135#_c_315_n N_VGND_c_1182_n 0.00376194f $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_416 N_A_154_135#_c_304_n N_VGND_c_1134_n 0.00467453f $X=4.24 $Y=1.35 $X2=0
+ $Y2=0
cc_417 N_A_154_135#_c_305_n N_VGND_c_1134_n 0.00405273f $X=4.67 $Y=1.35 $X2=0
+ $Y2=0
cc_418 N_A_154_135#_c_302_n N_VGND_c_1137_n 0.00505379f $X=3.38 $Y=1.35 $X2=0
+ $Y2=0
cc_419 N_A_154_135#_c_303_n N_VGND_c_1137_n 0.00505379f $X=3.81 $Y=1.35 $X2=0
+ $Y2=0
cc_420 N_A_154_135#_c_304_n N_VGND_c_1137_n 0.00505379f $X=4.24 $Y=1.35 $X2=0
+ $Y2=0
cc_421 N_A_154_135#_c_305_n N_VGND_c_1137_n 0.00424518f $X=4.67 $Y=1.35 $X2=0
+ $Y2=0
cc_422 N_A_154_135#_c_309_n N_VGND_c_1137_n 0.0103323f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_423 N_A_154_135#_c_311_n N_A_1346_123#_c_1261_n 0.0672585f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_424 N_A_154_135#_c_380_p N_A_1346_123#_c_1261_n 0.0136942f $X=8.28 $Y=0.76
+ $X2=0 $Y2=0
cc_425 N_A_154_135#_c_310_n N_A_1346_123#_c_1262_n 0.00406848f $X=6.005 $Y=1.6
+ $X2=0 $Y2=0
cc_426 N_A_154_135#_c_311_n N_A_1346_123#_c_1262_n 0.0273383f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_427 N_A_154_135#_c_314_n N_A_1346_123#_c_1262_n 6.69459e-19 $X=5.85 $Y=1.215
+ $X2=0 $Y2=0
cc_428 N_A_154_135#_c_380_p N_A_1346_123#_c_1263_n 0.0329533f $X=8.28 $Y=0.76
+ $X2=0 $Y2=0
cc_429 N_A_154_135#_M1011_d N_A_1346_123#_c_1264_n 0.00176461f $X=8.14 $Y=0.38
+ $X2=0 $Y2=0
cc_430 N_A_154_135#_c_380_p N_A_1346_123#_c_1264_n 0.0159805f $X=8.28 $Y=0.76
+ $X2=0 $Y2=0
cc_431 N_A_154_135#_c_380_p N_A_1346_123#_c_1266_n 0.0166977f $X=8.28 $Y=0.76
+ $X2=0 $Y2=0
cc_432 N_C1_c_516_n N_B2_c_588_n 0.0346059f $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_433 N_C1_c_516_n N_B2_M1016_g 0.00456705f $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_434 N_C1_c_516_n N_B2_c_582_n 0.0125599f $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_435 N_C1_M1026_g N_B2_c_586_n 8.38383e-19 $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_436 N_C1_M1026_g N_B2_c_587_n 0.0107847f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_437 N_C1_c_517_n N_VPWR_c_737_n 0.00278271f $X=5.86 $Y=1.885 $X2=0 $Y2=0
cc_438 N_C1_c_516_n N_VPWR_c_737_n 0.00278271f $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_439 N_C1_c_517_n N_VPWR_c_723_n 0.00358624f $X=5.86 $Y=1.885 $X2=0 $Y2=0
cc_440 N_C1_c_516_n N_VPWR_c_723_n 0.00353907f $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_441 N_C1_c_517_n N_A_157_376#_c_812_n 0.0167984f $X=5.86 $Y=1.885 $X2=0 $Y2=0
cc_442 N_C1_c_515_n N_A_157_376#_c_812_n 0.00108599f $X=6.065 $Y=1.515 $X2=0
+ $Y2=0
cc_443 N_C1_c_516_n N_A_157_376#_c_812_n 0.0124639f $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_444 C1 N_A_157_376#_c_812_n 0.0227239f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_445 N_C1_c_516_n N_A_157_376#_c_813_n 5.0035e-19 $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_446 N_C1_c_516_n N_A_157_376#_c_836_n 0.00104f $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_447 C1 N_A_1102_392#_M1003_s 0.00470299f $X=5.435 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_448 N_C1_c_517_n N_A_1102_392#_c_1024_n 0.0151248f $X=5.86 $Y=1.885 $X2=0
+ $Y2=0
cc_449 N_C1_c_516_n N_A_1102_392#_c_1024_n 0.0142207f $X=6.31 $Y=1.885 $X2=0
+ $Y2=0
cc_450 N_C1_M1024_g N_VGND_c_1122_n 0.00563785f $X=5.56 $Y=0.92 $X2=0 $Y2=0
cc_451 N_C1_M1026_g N_VGND_c_1123_n 0.00379263f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_452 N_C1_M1026_g N_VGND_c_1124_n 0.00215221f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_453 N_C1_c_516_n N_VGND_c_1124_n 0.00291802f $X=6.31 $Y=1.885 $X2=0 $Y2=0
cc_454 N_C1_M1024_g N_VGND_c_1131_n 0.00412501f $X=5.56 $Y=0.92 $X2=0 $Y2=0
cc_455 N_C1_M1026_g N_VGND_c_1131_n 0.00412501f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_456 N_C1_M1026_g N_VGND_c_1182_n 0.00298414f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_457 N_C1_c_514_n N_VGND_c_1182_n 0.0031599f $X=6.22 $Y=1.515 $X2=0 $Y2=0
cc_458 N_C1_M1024_g N_VGND_c_1137_n 0.00476395f $X=5.56 $Y=0.92 $X2=0 $Y2=0
cc_459 N_C1_M1026_g N_VGND_c_1137_n 0.00476395f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_460 N_C1_M1026_g N_A_1346_123#_c_1262_n 3.77674e-19 $X=5.99 $Y=0.92 $X2=0
+ $Y2=0
cc_461 N_B2_c_590_n N_B1_c_678_n 0.0178961f $X=7.21 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_462 N_B2_c_577_n N_B1_M1011_g 0.0131785f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_463 N_B2_c_580_n N_B1_c_675_n 0.0115034f $X=7.475 $Y=1.625 $X2=0 $Y2=0
cc_464 N_B2_c_581_n N_B1_c_675_n 0.0131785f $X=7.575 $Y=1.33 $X2=0 $Y2=0
cc_465 N_B2_c_583_n N_B1_c_675_n 0.00304467f $X=7.21 $Y=1.755 $X2=0 $Y2=0
cc_466 N_B2_c_588_n N_VPWR_c_737_n 0.00278271f $X=6.76 $Y=1.885 $X2=0 $Y2=0
cc_467 N_B2_c_590_n N_VPWR_c_737_n 0.00278271f $X=7.21 $Y=1.885 $X2=0 $Y2=0
cc_468 N_B2_c_588_n N_VPWR_c_723_n 0.00353907f $X=6.76 $Y=1.885 $X2=0 $Y2=0
cc_469 N_B2_c_590_n N_VPWR_c_723_n 0.00355937f $X=7.21 $Y=1.885 $X2=0 $Y2=0
cc_470 N_B2_c_588_n N_A_157_376#_c_812_n 0.0105104f $X=6.76 $Y=1.885 $X2=0 $Y2=0
cc_471 N_B2_c_588_n N_A_157_376#_c_813_n 0.00344562f $X=6.76 $Y=1.885 $X2=0
+ $Y2=0
cc_472 N_B2_c_578_n N_A_157_376#_c_813_n 0.00619098f $X=7.01 $Y=1.7 $X2=0 $Y2=0
cc_473 N_B2_c_590_n N_A_157_376#_c_813_n 6.83942e-19 $X=7.21 $Y=1.885 $X2=0
+ $Y2=0
cc_474 N_B2_c_582_n N_A_157_376#_c_813_n 3.81424e-19 $X=6.76 $Y=1.7 $X2=0 $Y2=0
cc_475 N_B2_c_583_n N_A_157_376#_c_813_n 4.69291e-19 $X=7.21 $Y=1.755 $X2=0
+ $Y2=0
cc_476 N_B2_c_588_n N_A_157_376#_c_836_n 0.00514748f $X=6.76 $Y=1.885 $X2=0
+ $Y2=0
cc_477 N_B2_c_590_n N_A_157_376#_c_836_n 0.0089426f $X=7.21 $Y=1.885 $X2=0 $Y2=0
cc_478 N_B2_c_590_n N_A_157_376#_c_814_n 0.0130998f $X=7.21 $Y=1.885 $X2=0 $Y2=0
cc_479 N_B2_c_583_n N_A_157_376#_c_814_n 0.0066701f $X=7.21 $Y=1.755 $X2=0 $Y2=0
cc_480 N_B2_c_588_n N_A_157_376#_c_856_n 7.24124e-19 $X=6.76 $Y=1.885 $X2=0
+ $Y2=0
cc_481 N_B2_c_590_n N_A_157_376#_c_856_n 0.0051685f $X=7.21 $Y=1.885 $X2=0 $Y2=0
cc_482 N_B2_c_588_n N_A_1102_392#_c_1025_n 0.00774277f $X=6.76 $Y=1.885 $X2=0
+ $Y2=0
cc_483 N_B2_c_590_n N_A_1102_392#_c_1025_n 0.0146423f $X=7.21 $Y=1.885 $X2=0
+ $Y2=0
cc_484 N_B2_c_590_n N_A_1102_392#_c_1036_n 0.00957545f $X=7.21 $Y=1.885 $X2=0
+ $Y2=0
cc_485 N_B2_c_588_n N_A_1102_392#_c_1028_n 0.0055162f $X=6.76 $Y=1.885 $X2=0
+ $Y2=0
cc_486 N_B2_c_590_n N_A_1102_392#_c_1028_n 7.34383e-19 $X=7.21 $Y=1.885 $X2=0
+ $Y2=0
cc_487 N_B2_c_585_n N_VGND_c_1123_n 0.0243585f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_488 N_B2_c_586_n N_VGND_c_1123_n 0.00566684f $X=6.635 $Y=0.2 $X2=0 $Y2=0
cc_489 N_B2_c_587_n N_VGND_c_1123_n 0.00167326f $X=6.635 $Y=0.505 $X2=0 $Y2=0
cc_490 N_B2_c_587_n N_VGND_c_1124_n 2.51918e-19 $X=6.635 $Y=0.505 $X2=0 $Y2=0
cc_491 N_B2_c_577_n N_VGND_c_1125_n 0.0193089f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_492 N_B2_M1016_g N_VGND_c_1125_n 0.00161245f $X=7.085 $Y=0.935 $X2=0 $Y2=0
cc_493 N_B2_c_581_n N_VGND_c_1125_n 0.00832159f $X=7.575 $Y=1.33 $X2=0 $Y2=0
cc_494 N_B2_c_584_n N_VGND_c_1125_n 4.2102e-19 $X=7.575 $Y=1.405 $X2=0 $Y2=0
cc_495 N_B2_c_585_n N_VGND_c_1125_n 0.029476f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_496 N_B2_c_585_n N_VGND_c_1182_n 0.00386879f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_497 N_B2_c_586_n N_VGND_c_1182_n 0.00127982f $X=6.635 $Y=0.2 $X2=0 $Y2=0
cc_498 N_B2_c_585_n N_VGND_c_1135_n 0.0366677f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_499 N_B2_c_586_n N_VGND_c_1135_n 0.0181591f $X=6.635 $Y=0.2 $X2=0 $Y2=0
cc_500 N_B2_c_577_n N_VGND_c_1136_n 0.00693208f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_501 N_B2_c_577_n N_VGND_c_1137_n 0.0256169f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_502 N_B2_M1016_g N_VGND_c_1137_n 7.07849e-19 $X=7.085 $Y=0.935 $X2=0 $Y2=0
cc_503 N_B2_c_585_n N_VGND_c_1137_n 0.0191717f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_504 N_B2_c_586_n N_VGND_c_1137_n 0.0100038f $X=6.635 $Y=0.2 $X2=0 $Y2=0
cc_505 N_B2_c_585_n N_A_1346_123#_M1014_d 0.00190525f $X=6.845 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_506 N_B2_c_577_n N_A_1346_123#_c_1278_n 3.49074e-19 $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_507 N_B2_M1016_g N_A_1346_123#_c_1278_n 0.00657116f $X=7.085 $Y=0.935 $X2=0
+ $Y2=0
cc_508 N_B2_c_581_n N_A_1346_123#_c_1278_n 5.93148e-19 $X=7.575 $Y=1.33 $X2=0
+ $Y2=0
cc_509 N_B2_c_585_n N_A_1346_123#_c_1278_n 0.0156219f $X=6.845 $Y=0.38 $X2=0
+ $Y2=0
cc_510 N_B2_c_586_n N_A_1346_123#_c_1278_n 0.00127917f $X=6.635 $Y=0.2 $X2=0
+ $Y2=0
cc_511 N_B2_c_587_n N_A_1346_123#_c_1278_n 0.00526654f $X=6.635 $Y=0.505 $X2=0
+ $Y2=0
cc_512 N_B2_M1016_g N_A_1346_123#_c_1261_n 0.0109993f $X=7.085 $Y=0.935 $X2=0
+ $Y2=0
cc_513 N_B2_c_581_n N_A_1346_123#_c_1261_n 0.00932666f $X=7.575 $Y=1.33 $X2=0
+ $Y2=0
cc_514 N_B2_c_583_n N_A_1346_123#_c_1261_n 3.92729e-19 $X=7.21 $Y=1.755 $X2=0
+ $Y2=0
cc_515 N_B2_c_584_n N_A_1346_123#_c_1261_n 0.00873336f $X=7.575 $Y=1.405 $X2=0
+ $Y2=0
cc_516 N_B2_c_585_n N_A_1346_123#_c_1261_n 2.22629e-19 $X=6.845 $Y=0.38 $X2=0
+ $Y2=0
cc_517 N_B2_M1016_g N_A_1346_123#_c_1262_n 0.00314813f $X=7.085 $Y=0.935 $X2=0
+ $Y2=0
cc_518 N_B2_c_582_n N_A_1346_123#_c_1262_n 0.00212048f $X=6.76 $Y=1.7 $X2=0
+ $Y2=0
cc_519 N_B2_c_587_n N_A_1346_123#_c_1262_n 0.00390184f $X=6.635 $Y=0.505 $X2=0
+ $Y2=0
cc_520 N_B2_c_581_n N_A_1346_123#_c_1263_n 0.0086474f $X=7.575 $Y=1.33 $X2=0
+ $Y2=0
cc_521 N_B2_c_577_n N_A_1346_123#_c_1265_n 0.0017897f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_522 N_B1_c_678_n N_VPWR_c_737_n 0.00278271f $X=7.95 $Y=1.885 $X2=0 $Y2=0
cc_523 N_B1_c_679_n N_VPWR_c_737_n 0.00278271f $X=8.44 $Y=1.885 $X2=0 $Y2=0
cc_524 N_B1_c_678_n N_VPWR_c_723_n 0.00356309f $X=7.95 $Y=1.885 $X2=0 $Y2=0
cc_525 N_B1_c_679_n N_VPWR_c_723_n 0.00358997f $X=8.44 $Y=1.885 $X2=0 $Y2=0
cc_526 N_B1_c_678_n N_A_157_376#_c_814_n 0.0130998f $X=7.95 $Y=1.885 $X2=0 $Y2=0
cc_527 N_B1_c_675_n N_A_157_376#_c_814_n 3.81992e-19 $X=8.57 $Y=1.51 $X2=0 $Y2=0
cc_528 N_B1_c_678_n N_A_157_376#_c_817_n 0.0154053f $X=7.95 $Y=1.885 $X2=0 $Y2=0
cc_529 N_B1_c_679_n N_A_157_376#_c_817_n 0.0108953f $X=8.44 $Y=1.885 $X2=0 $Y2=0
cc_530 N_B1_c_675_n N_A_157_376#_c_817_n 0.00308717f $X=8.57 $Y=1.51 $X2=0 $Y2=0
cc_531 N_B1_c_678_n N_A_1102_392#_c_1036_n 0.00976577f $X=7.95 $Y=1.885 $X2=0
+ $Y2=0
cc_532 N_B1_c_678_n N_A_1102_392#_c_1026_n 0.0148944f $X=7.95 $Y=1.885 $X2=0
+ $Y2=0
cc_533 N_B1_c_679_n N_A_1102_392#_c_1026_n 0.0139261f $X=8.44 $Y=1.885 $X2=0
+ $Y2=0
cc_534 N_B1_c_679_n N_A_1102_392#_c_1027_n 0.00670792f $X=8.44 $Y=1.885 $X2=0
+ $Y2=0
cc_535 N_B1_c_677_n N_A_1102_392#_c_1027_n 0.00301248f $X=9.115 $Y=1.465 $X2=0
+ $Y2=0
cc_536 N_B1_c_683_n N_A_1102_392#_c_1027_n 0.0178913f $X=9.095 $Y=1.48 $X2=0
+ $Y2=0
cc_537 N_B1_M1011_g N_VGND_c_1136_n 0.00390708f $X=8.065 $Y=0.7 $X2=0 $Y2=0
cc_538 N_B1_M1018_g N_VGND_c_1136_n 0.00390708f $X=8.495 $Y=0.7 $X2=0 $Y2=0
cc_539 N_B1_M1011_g N_VGND_c_1137_n 0.00542671f $X=8.065 $Y=0.7 $X2=0 $Y2=0
cc_540 N_B1_M1018_g N_VGND_c_1137_n 0.00542671f $X=8.495 $Y=0.7 $X2=0 $Y2=0
cc_541 N_B1_M1011_g N_A_1346_123#_c_1261_n 0.00164273f $X=8.065 $Y=0.7 $X2=0
+ $Y2=0
cc_542 N_B1_c_675_n N_A_1346_123#_c_1261_n 0.0020527f $X=8.57 $Y=1.51 $X2=0
+ $Y2=0
cc_543 N_B1_M1011_g N_A_1346_123#_c_1263_n 0.00195727f $X=8.065 $Y=0.7 $X2=0
+ $Y2=0
cc_544 N_B1_M1011_g N_A_1346_123#_c_1264_n 0.0123852f $X=8.065 $Y=0.7 $X2=0
+ $Y2=0
cc_545 N_B1_M1018_g N_A_1346_123#_c_1264_n 0.0135055f $X=8.495 $Y=0.7 $X2=0
+ $Y2=0
cc_546 N_B1_M1018_g N_A_1346_123#_c_1266_n 4.46492e-19 $X=8.495 $Y=0.7 $X2=0
+ $Y2=0
cc_547 N_B1_c_677_n N_A_1346_123#_c_1266_n 0.00691526f $X=9.115 $Y=1.465 $X2=0
+ $Y2=0
cc_548 N_B1_c_683_n N_A_1346_123#_c_1266_n 0.0186971f $X=9.095 $Y=1.48 $X2=0
+ $Y2=0
cc_549 N_VPWR_M1004_s N_A_157_376#_c_818_n 0.0170117f $X=1.355 $Y=1.88 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_739_n N_A_157_376#_c_818_n 0.0513372f $X=1.9 $Y=2.71 $X2=0 $Y2=0
cc_551 N_VPWR_M1015_s N_A_157_376#_c_812_n 0.00926123f $X=2.7 $Y=1.88 $X2=0
+ $Y2=0
cc_552 N_VPWR_M1017_d N_A_157_376#_c_812_n 0.00378605f $X=3.76 $Y=1.84 $X2=0
+ $Y2=0
cc_553 N_VPWR_M1025_d N_A_157_376#_c_812_n 0.00854919f $X=4.66 $Y=1.84 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_725_n N_A_157_376#_c_812_n 0.0214637f $X=3.01 $Y=2.8 $X2=0 $Y2=0
cc_555 N_VPWR_c_726_n N_A_157_376#_c_812_n 0.0168121f $X=3.91 $Y=2.8 $X2=0 $Y2=0
cc_556 N_VPWR_c_727_n N_A_157_376#_c_812_n 0.0215824f $X=4.81 $Y=2.8 $X2=0 $Y2=0
cc_557 N_VPWR_c_723_n N_A_157_376#_c_812_n 0.0697223f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_724_n N_A_157_376#_c_815_n 0.0387673f $X=0.485 $Y=2.345 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_736_n N_A_157_376#_c_815_n 0.0109716f $X=1.395 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_723_n N_A_157_376#_c_815_n 0.0114726f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_739_n N_A_157_376#_c_815_n 0.0118598f $X=1.9 $Y=2.71 $X2=0 $Y2=0
cc_562 N_VPWR_c_725_n N_A_157_376#_c_816_n 0.0106233f $X=3.01 $Y=2.8 $X2=0 $Y2=0
cc_563 N_VPWR_c_730_n N_A_157_376#_c_816_n 0.0109344f $X=2.845 $Y=3.33 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_723_n N_A_157_376#_c_816_n 0.0114592f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_739_n N_A_157_376#_c_816_n 0.0121364f $X=1.9 $Y=2.71 $X2=0 $Y2=0
cc_566 N_VPWR_c_724_n N_X_c_910_n 0.00313887f $X=0.485 $Y=2.345 $X2=0 $Y2=0
cc_567 N_VPWR_M1015_s N_X_c_922_n 0.00807578f $X=2.7 $Y=1.88 $X2=0 $Y2=0
cc_568 N_VPWR_M1017_d N_X_c_934_n 0.00362442f $X=3.76 $Y=1.84 $X2=0 $Y2=0
cc_569 N_VPWR_M1001_s N_X_c_912_n 0.00741318f $X=0.36 $Y=1.88 $X2=0 $Y2=0
cc_570 N_VPWR_M1004_s N_X_c_912_n 0.0169013f $X=1.355 $Y=1.88 $X2=0 $Y2=0
cc_571 N_VPWR_M1015_s N_X_c_912_n 0.00202056f $X=2.7 $Y=1.88 $X2=0 $Y2=0
cc_572 N_VPWR_c_724_n N_X_c_912_n 0.019145f $X=0.485 $Y=2.345 $X2=0 $Y2=0
cc_573 N_VPWR_c_727_n N_A_1102_392#_c_1024_n 0.0157109f $X=4.81 $Y=2.8 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_737_n N_A_1102_392#_c_1024_n 0.128567f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_723_n N_A_1102_392#_c_1024_n 0.0715883f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_737_n N_A_1102_392#_c_1026_n 0.0701352f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_723_n N_A_1102_392#_c_1026_n 0.0393644f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_737_n N_A_1102_392#_c_1029_n 0.0236566f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_723_n N_A_1102_392#_c_1029_n 0.0128296f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_580 N_A_157_376#_c_812_n N_X_M1000_s 0.00545306f $X=6.82 $Y=2.445 $X2=0 $Y2=0
cc_581 N_A_157_376#_c_812_n N_X_M1019_s 0.00545306f $X=6.82 $Y=2.445 $X2=0 $Y2=0
cc_582 N_A_157_376#_c_812_n N_X_c_922_n 0.0935511f $X=6.82 $Y=2.445 $X2=0 $Y2=0
cc_583 N_A_157_376#_M1001_d N_X_c_912_n 0.00815711f $X=0.785 $Y=1.88 $X2=0 $Y2=0
cc_584 N_A_157_376#_M1013_d N_X_c_912_n 0.00380424f $X=2.25 $Y=1.88 $X2=0 $Y2=0
cc_585 N_A_157_376#_c_818_n N_X_c_912_n 0.0640645f $X=2.235 $Y=2.345 $X2=0 $Y2=0
cc_586 N_A_157_376#_c_812_n N_X_c_912_n 0.0110789f $X=6.82 $Y=2.445 $X2=0 $Y2=0
cc_587 N_A_157_376#_c_815_n N_X_c_912_n 0.0219827f $X=1.055 $Y=2.345 $X2=0 $Y2=0
cc_588 N_A_157_376#_c_816_n N_X_c_912_n 0.0172489f $X=2.4 $Y=2.345 $X2=0 $Y2=0
cc_589 N_A_157_376#_c_812_n N_A_1102_392#_M1003_s 0.00545233f $X=6.82 $Y=2.445
+ $X2=-0.19 $Y2=1.66
cc_590 N_A_157_376#_c_812_n N_A_1102_392#_M1006_s 0.00561849f $X=6.82 $Y=2.445
+ $X2=0 $Y2=0
cc_591 N_A_157_376#_c_814_n N_A_1102_392#_M1009_s 0.0110306f $X=8.01 $Y=2.025
+ $X2=0 $Y2=0
cc_592 N_A_157_376#_c_812_n N_A_1102_392#_c_1024_n 0.0693779f $X=6.82 $Y=2.445
+ $X2=0 $Y2=0
cc_593 N_A_157_376#_M1008_d N_A_1102_392#_c_1025_n 0.00197722f $X=6.835 $Y=1.96
+ $X2=0 $Y2=0
cc_594 N_A_157_376#_c_812_n N_A_1102_392#_c_1025_n 0.00368894f $X=6.82 $Y=2.445
+ $X2=0 $Y2=0
cc_595 N_A_157_376#_c_856_n N_A_1102_392#_c_1025_n 0.0156803f $X=6.985 $Y=2.445
+ $X2=0 $Y2=0
cc_596 N_A_157_376#_c_836_n N_A_1102_392#_c_1036_n 0.00426962f $X=6.985 $Y=2.36
+ $X2=0 $Y2=0
cc_597 N_A_157_376#_c_814_n N_A_1102_392#_c_1036_n 0.0266856f $X=8.01 $Y=2.025
+ $X2=0 $Y2=0
cc_598 N_A_157_376#_c_856_n N_A_1102_392#_c_1036_n 0.020576f $X=6.985 $Y=2.445
+ $X2=0 $Y2=0
cc_599 N_A_157_376#_c_817_n N_A_1102_392#_c_1036_n 0.0260984f $X=8.195 $Y=2.105
+ $X2=0 $Y2=0
cc_600 N_A_157_376#_M1010_d N_A_1102_392#_c_1026_n 0.00240242f $X=8.025 $Y=1.96
+ $X2=0 $Y2=0
cc_601 N_A_157_376#_c_817_n N_A_1102_392#_c_1026_n 0.0191222f $X=8.195 $Y=2.105
+ $X2=0 $Y2=0
cc_602 N_A_157_376#_c_817_n N_A_1102_392#_c_1027_n 0.0543691f $X=8.195 $Y=2.105
+ $X2=0 $Y2=0
cc_603 N_X_c_905_n N_A_71_135#_M1005_s 0.0019963f $X=2.975 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_604 N_X_c_906_n N_A_71_135#_M1005_s 7.27654e-19 $X=0.385 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_605 N_X_c_905_n N_A_71_135#_M1007_s 0.00206067f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_606 N_X_c_905_n N_A_71_135#_M1022_d 0.00201585f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_607 N_X_c_905_n N_A_71_135#_c_1069_n 0.012018f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_608 N_X_c_905_n N_A_71_135#_c_1074_n 0.00908056f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_609 N_X_c_905_n N_A_71_135#_c_1066_n 0.0443333f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_610 X N_A_71_135#_c_1066_n 0.00129662f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_611 N_X_c_909_n N_A_71_135#_c_1066_n 0.00793711f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_612 N_X_c_905_n N_A_71_135#_c_1067_n 0.00564678f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_613 N_X_c_905_n N_A_71_135#_c_1085_n 0.00591085f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_614 X N_A_71_135#_c_1085_n 0.00128755f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_615 N_X_c_909_n N_A_71_135#_c_1085_n 9.21622e-19 $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_616 N_X_c_905_n N_A_71_135#_c_1068_n 0.00835176f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_617 N_X_c_906_n N_A_71_135#_c_1068_n 0.00187568f $X=0.385 $Y=1.295 $X2=0
+ $Y2=0
cc_618 N_X_c_907_n N_A_71_135#_c_1068_n 0.0027311f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_619 N_X_c_905_n N_VGND_M1022_s 0.00372485f $X=2.975 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_620 N_X_c_940_n N_VGND_M1027_s 6.98766e-19 $X=3.43 $Y=1.095 $X2=0 $Y2=0
cc_621 N_X_c_905_n N_VGND_M1027_s 3.42314e-19 $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_622 X N_VGND_M1027_s 0.00254293f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_623 N_X_c_909_n N_VGND_M1027_s 0.00512514f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_624 N_X_c_946_n N_VGND_M1012_s 0.00330483f $X=4.29 $Y=1.095 $X2=0 $Y2=0
cc_625 N_X_c_940_n N_VGND_c_1120_n 9.87298e-19 $X=3.43 $Y=1.095 $X2=0 $Y2=0
cc_626 N_X_c_903_n N_VGND_c_1120_n 0.0165971f $X=3.595 $Y=0.645 $X2=0 $Y2=0
cc_627 X N_VGND_c_1120_n 0.00158234f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_628 N_X_c_909_n N_VGND_c_1120_n 0.0172527f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_629 N_X_c_903_n N_VGND_c_1121_n 0.0164685f $X=3.595 $Y=0.645 $X2=0 $Y2=0
cc_630 N_X_c_946_n N_VGND_c_1121_n 0.0135055f $X=4.29 $Y=1.095 $X2=0 $Y2=0
cc_631 N_X_c_904_n N_VGND_c_1121_n 0.013052f $X=4.455 $Y=0.645 $X2=0 $Y2=0
cc_632 N_X_c_904_n N_VGND_c_1122_n 0.0201101f $X=4.455 $Y=0.645 $X2=0 $Y2=0
cc_633 N_X_c_905_n N_VGND_c_1128_n 0.0103398f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_634 N_X_c_903_n N_VGND_c_1129_n 0.0105983f $X=3.595 $Y=0.645 $X2=0 $Y2=0
cc_635 N_X_c_904_n N_VGND_c_1134_n 0.00718756f $X=4.455 $Y=0.645 $X2=0 $Y2=0
cc_636 N_X_c_903_n N_VGND_c_1137_n 0.0113894f $X=3.595 $Y=0.645 $X2=0 $Y2=0
cc_637 N_X_c_904_n N_VGND_c_1137_n 0.0083989f $X=4.455 $Y=0.645 $X2=0 $Y2=0
cc_638 N_A_71_135#_c_1066_n N_VGND_M1022_s 9.8611e-19 $X=2.51 $Y=1.325 $X2=-0.19
+ $Y2=-0.245
cc_639 N_A_71_135#_c_1069_n N_VGND_c_1126_n 0.0105986f $X=1.255 $Y=0.82 $X2=0
+ $Y2=0
cc_640 N_A_71_135#_c_1068_n N_VGND_c_1126_n 0.00458739f $X=0.48 $Y=0.83 $X2=0
+ $Y2=0
cc_641 N_A_71_135#_c_1074_n N_VGND_c_1128_n 0.00104849f $X=1.34 $Y=1.035 $X2=0
+ $Y2=0
cc_642 N_A_71_135#_c_1066_n N_VGND_c_1128_n 0.0269989f $X=2.51 $Y=1.325 $X2=0
+ $Y2=0
cc_643 N_A_71_135#_c_1069_n N_VGND_c_1137_n 0.0226601f $X=1.255 $Y=0.82 $X2=0
+ $Y2=0
cc_644 N_A_71_135#_c_1085_n N_VGND_c_1137_n 5.77272e-19 $X=2.675 $Y=1.055 $X2=0
+ $Y2=0
cc_645 N_A_71_135#_c_1068_n N_VGND_c_1137_n 0.00719958f $X=0.48 $Y=0.83 $X2=0
+ $Y2=0
cc_646 N_VGND_c_1124_n N_A_1346_123#_c_1278_n 0.0108698f $X=6.44 $Y=1.115 $X2=0
+ $Y2=0
cc_647 N_VGND_c_1137_n N_A_1346_123#_c_1278_n 8.15299e-19 $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_648 N_VGND_c_1125_n N_A_1346_123#_c_1261_n 0.0205307f $X=7.3 $Y=0.925 $X2=0
+ $Y2=0
cc_649 N_VGND_c_1124_n N_A_1346_123#_c_1262_n 0.00157382f $X=6.44 $Y=1.115 $X2=0
+ $Y2=0
cc_650 N_VGND_c_1125_n N_A_1346_123#_c_1263_n 0.0442411f $X=7.3 $Y=0.925 $X2=0
+ $Y2=0
cc_651 N_VGND_c_1136_n N_A_1346_123#_c_1264_n 0.0650231f $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_652 N_VGND_c_1137_n N_A_1346_123#_c_1264_n 0.037428f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_653 N_VGND_c_1125_n N_A_1346_123#_c_1265_n 0.0122034f $X=7.3 $Y=0.925 $X2=0
+ $Y2=0
cc_654 N_VGND_c_1136_n N_A_1346_123#_c_1265_n 0.0179217f $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_655 N_VGND_c_1137_n N_A_1346_123#_c_1265_n 0.00971942f $X=9.36 $Y=0 $X2=0
+ $Y2=0
