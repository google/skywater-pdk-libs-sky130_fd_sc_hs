* File: sky130_fd_sc_hs__nand3b_1.pxi.spice
* Created: Thu Aug 27 20:51:17 2020
* 
x_PM_SKY130_FD_SC_HS__NAND3B_1%A_N N_A_N_M1003_g N_A_N_c_48_n N_A_N_M1005_g A_N
+ N_A_N_c_49_n PM_SKY130_FD_SC_HS__NAND3B_1%A_N
x_PM_SKY130_FD_SC_HS__NAND3B_1%C N_C_c_73_n N_C_M1002_g N_C_M1006_g C N_C_c_75_n
+ PM_SKY130_FD_SC_HS__NAND3B_1%C
x_PM_SKY130_FD_SC_HS__NAND3B_1%B N_B_M1007_g N_B_c_102_n N_B_M1004_g B
+ N_B_c_103_n PM_SKY130_FD_SC_HS__NAND3B_1%B
x_PM_SKY130_FD_SC_HS__NAND3B_1%A_27_116# N_A_27_116#_M1003_s N_A_27_116#_M1005_s
+ N_A_27_116#_M1000_g N_A_27_116#_c_135_n N_A_27_116#_M1001_g
+ N_A_27_116#_c_136_n N_A_27_116#_c_137_n N_A_27_116#_c_138_n
+ N_A_27_116#_c_139_n N_A_27_116#_c_143_n N_A_27_116#_c_140_n
+ N_A_27_116#_c_141_n PM_SKY130_FD_SC_HS__NAND3B_1%A_27_116#
x_PM_SKY130_FD_SC_HS__NAND3B_1%VPWR N_VPWR_M1005_d N_VPWR_M1004_d N_VPWR_c_197_n
+ N_VPWR_c_198_n N_VPWR_c_199_n N_VPWR_c_200_n N_VPWR_c_201_n N_VPWR_c_202_n
+ VPWR N_VPWR_c_203_n N_VPWR_c_196_n PM_SKY130_FD_SC_HS__NAND3B_1%VPWR
x_PM_SKY130_FD_SC_HS__NAND3B_1%Y N_Y_M1000_d N_Y_M1002_d N_Y_M1001_d N_Y_c_237_n
+ N_Y_c_233_n N_Y_c_243_n N_Y_c_231_n Y Y Y N_Y_c_235_n N_Y_c_232_n
+ PM_SKY130_FD_SC_HS__NAND3B_1%Y
x_PM_SKY130_FD_SC_HS__NAND3B_1%VGND N_VGND_M1003_d N_VGND_c_272_n VGND
+ N_VGND_c_273_n N_VGND_c_274_n N_VGND_c_275_n N_VGND_c_276_n
+ PM_SKY130_FD_SC_HS__NAND3B_1%VGND
cc_1 VNB N_A_N_M1003_g 0.0310639f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.855
cc_2 VNB N_A_N_c_48_n 0.0285737f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.765
cc_3 VNB N_A_N_c_49_n 0.00453475f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_4 VNB N_C_c_73_n 0.0270203f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_5 VNB N_C_M1006_g 0.0255815f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.26
cc_6 VNB N_C_c_75_n 0.00176544f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_7 VNB N_B_M1007_g 0.0233178f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.855
cc_8 VNB N_B_c_102_n 0.0247044f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.765
cc_9 VNB N_B_c_103_n 0.00404949f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_10 VNB N_A_27_116#_M1000_g 0.0267595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_116#_c_135_n 0.0343849f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_12 VNB N_A_27_116#_c_136_n 0.0191713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_116#_c_137_n 0.0257611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_116#_c_138_n 0.00199818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_116#_c_139_n 0.0111529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_116#_c_140_n 0.0238989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_116#_c_141_n 0.00579502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_196_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_231_n 0.03984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_232_n 0.0239082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_272_n 0.0174336f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.26
cc_22 VNB N_VGND_c_273_n 0.0181018f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.515
cc_23 VNB N_VGND_c_274_n 0.0508477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_275_n 0.21221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_276_n 0.0129456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_A_N_c_48_n 0.0332688f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.765
cc_27 VPB N_A_N_c_49_n 0.00601631f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_28 VPB N_C_c_73_n 0.0274529f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_29 VPB N_C_c_75_n 0.00404813f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_30 VPB N_B_c_102_n 0.0272948f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.765
cc_31 VPB N_B_c_103_n 0.00376788f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_32 VPB N_A_27_116#_c_135_n 0.0291369f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_33 VPB N_A_27_116#_c_143_n 0.0414281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_27_116#_c_140_n 0.0140293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_197_n 0.0195801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_198_n 0.00900305f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_37 VPB N_VPWR_c_199_n 0.0255433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_200_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_201_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_202_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_203_n 0.0220385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_196_n 0.0650812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_Y_c_233_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_44 VPB Y 0.0434383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_Y_c_235_n 0.0171662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_232_n 0.00787282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 N_A_N_c_48_n N_C_c_73_n 0.0413213f $X=0.66 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_48 N_A_N_c_49_n N_C_c_73_n 0.00231967f $X=0.61 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_49 N_A_N_M1003_g N_C_M1006_g 0.00972195f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_50 N_A_N_c_48_n N_C_c_75_n 6.90406e-19 $X=0.66 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A_N_c_49_n N_C_c_75_n 0.0334549f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_52 N_A_N_M1003_g N_A_27_116#_c_136_n 0.00199671f $X=0.495 $Y=0.855 $X2=0
+ $Y2=0
cc_53 N_A_N_M1003_g N_A_27_116#_c_137_n 0.0161994f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_54 N_A_N_c_48_n N_A_27_116#_c_137_n 0.0013821f $X=0.66 $Y=1.765 $X2=0 $Y2=0
cc_55 N_A_N_c_49_n N_A_27_116#_c_137_n 0.0262311f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_56 N_A_N_c_48_n N_A_27_116#_c_143_n 0.011153f $X=0.66 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A_N_c_49_n N_A_27_116#_c_143_n 0.0108778f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_58 N_A_N_M1003_g N_A_27_116#_c_140_n 0.0129934f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_59 N_A_N_c_48_n N_A_27_116#_c_140_n 0.00405327f $X=0.66 $Y=1.765 $X2=0 $Y2=0
cc_60 N_A_N_c_49_n N_A_27_116#_c_140_n 0.0331559f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_61 N_A_N_c_48_n N_VPWR_c_197_n 0.0103799f $X=0.66 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A_N_c_49_n N_VPWR_c_197_n 0.00248668f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_63 N_A_N_c_48_n N_VPWR_c_199_n 0.00393873f $X=0.66 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_N_c_48_n N_VPWR_c_196_n 0.00462577f $X=0.66 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A_N_M1003_g N_VGND_c_272_n 0.0112592f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_66 N_A_N_M1003_g N_VGND_c_273_n 0.00365567f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_67 N_A_N_M1003_g N_VGND_c_275_n 0.00404919f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_68 N_C_M1006_g N_B_M1007_g 0.0388863f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_69 N_C_c_73_n N_B_c_102_n 0.0552437f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_70 N_C_c_75_n N_B_c_102_n 7.44632e-19 $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_71 N_C_c_73_n N_B_c_103_n 0.0023886f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_72 N_C_c_75_n N_B_c_103_n 0.028624f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_73 N_C_c_73_n N_A_27_116#_c_137_n 0.00121615f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_74 N_C_M1006_g N_A_27_116#_c_137_n 0.0155047f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_75 N_C_c_75_n N_A_27_116#_c_137_n 0.021788f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_76 N_C_c_73_n N_VPWR_c_197_n 0.0128569f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_77 N_C_c_75_n N_VPWR_c_197_n 0.00953283f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_78 N_C_c_73_n N_VPWR_c_201_n 0.00445602f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_79 N_C_c_73_n N_VPWR_c_196_n 0.00861803f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_80 N_C_c_73_n N_Y_c_237_n 0.00184961f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_81 N_C_c_75_n N_Y_c_237_n 0.00223417f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_82 N_C_c_73_n N_Y_c_233_n 0.00871372f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_83 N_C_M1006_g N_VGND_c_272_n 0.01739f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_84 N_C_M1006_g N_VGND_c_274_n 0.00468165f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_85 N_C_M1006_g N_VGND_c_275_n 0.00453141f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_86 N_B_M1007_g N_A_27_116#_M1000_g 0.0344152f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_87 N_B_c_102_n N_A_27_116#_c_135_n 0.0544801f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_88 N_B_c_103_n N_A_27_116#_c_135_n 0.00282136f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_89 N_B_M1007_g N_A_27_116#_c_137_n 0.0154731f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_90 N_B_c_102_n N_A_27_116#_c_137_n 0.00121529f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_91 N_B_c_103_n N_A_27_116#_c_137_n 0.0232305f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_92 N_B_M1007_g N_A_27_116#_c_138_n 0.00296442f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_93 N_B_M1007_g N_A_27_116#_c_141_n 5.87559e-19 $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_94 N_B_c_102_n N_A_27_116#_c_141_n 0.00170526f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_95 N_B_c_103_n N_A_27_116#_c_141_n 0.0240984f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_96 N_B_c_102_n N_VPWR_c_198_n 0.00598632f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B_c_102_n N_VPWR_c_201_n 0.00445602f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_98 N_B_c_102_n N_VPWR_c_196_n 0.00857909f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B_c_102_n N_Y_c_237_n 4.2644e-19 $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_100 N_B_c_103_n N_Y_c_237_n 0.00354605f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_101 N_B_c_102_n N_Y_c_233_n 0.010308f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_102 N_B_c_102_n N_Y_c_243_n 0.0130725f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_103 N_B_c_103_n N_Y_c_243_n 0.0193106f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_104 N_B_M1007_g N_Y_c_231_n 0.00193784f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_105 N_B_c_102_n N_Y_c_235_n 0.00133299f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_106 N_B_M1007_g N_VGND_c_272_n 0.00269744f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_107 N_B_M1007_g N_VGND_c_274_n 0.00563421f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_108 N_B_M1007_g N_VGND_c_275_n 0.00539454f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_109 N_A_27_116#_c_143_n N_VPWR_c_197_n 0.0519547f $X=0.435 $Y=2.115 $X2=0
+ $Y2=0
cc_110 N_A_27_116#_c_135_n N_VPWR_c_198_n 0.00737447f $X=2.245 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_27_116#_c_143_n N_VPWR_c_199_n 0.0100559f $X=0.435 $Y=2.115 $X2=0
+ $Y2=0
cc_112 N_A_27_116#_c_135_n N_VPWR_c_203_n 0.00445602f $X=2.245 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A_27_116#_c_135_n N_VPWR_c_196_n 0.00861677f $X=2.245 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_27_116#_c_143_n N_VPWR_c_196_n 0.0149991f $X=0.435 $Y=2.115 $X2=0
+ $Y2=0
cc_115 N_A_27_116#_c_135_n N_Y_c_233_n 6.63528e-19 $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_27_116#_c_135_n N_Y_c_243_n 0.0137201f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_27_116#_c_141_n N_Y_c_243_n 0.00898653f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_118 N_A_27_116#_M1000_g N_Y_c_231_n 0.0222284f $X=2.2 $Y=0.76 $X2=0 $Y2=0
cc_119 N_A_27_116#_c_135_n N_Y_c_231_n 0.00328304f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_27_116#_c_137_n N_Y_c_231_n 0.0145858f $X=2.085 $Y=1.065 $X2=0 $Y2=0
cc_121 N_A_27_116#_c_141_n N_Y_c_231_n 0.00703632f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_122 N_A_27_116#_c_135_n Y 0.0116155f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_27_116#_c_135_n N_Y_c_235_n 0.00721634f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_27_116#_c_141_n N_Y_c_235_n 0.0125024f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_125 N_A_27_116#_M1000_g N_Y_c_232_n 0.00203887f $X=2.2 $Y=0.76 $X2=0 $Y2=0
cc_126 N_A_27_116#_c_135_n N_Y_c_232_n 0.00598143f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_27_116#_c_138_n N_Y_c_232_n 0.00479588f $X=2.17 $Y=1.32 $X2=0 $Y2=0
cc_128 N_A_27_116#_c_141_n N_Y_c_232_n 0.0249903f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_129 N_A_27_116#_c_137_n N_VGND_M1003_d 0.00761754f $X=2.085 $Y=1.065
+ $X2=-0.19 $Y2=-0.245
cc_130 N_A_27_116#_c_136_n N_VGND_c_272_n 0.0112316f $X=0.28 $Y=0.855 $X2=0
+ $Y2=0
cc_131 N_A_27_116#_c_137_n N_VGND_c_272_n 0.0451464f $X=2.085 $Y=1.065 $X2=0
+ $Y2=0
cc_132 N_A_27_116#_c_136_n N_VGND_c_273_n 0.00637154f $X=0.28 $Y=0.855 $X2=0
+ $Y2=0
cc_133 N_A_27_116#_M1000_g N_VGND_c_274_n 0.0053639f $X=2.2 $Y=0.76 $X2=0 $Y2=0
cc_134 N_A_27_116#_M1000_g N_VGND_c_275_n 0.00539454f $X=2.2 $Y=0.76 $X2=0 $Y2=0
cc_135 N_A_27_116#_c_136_n N_VGND_c_275_n 0.00857079f $X=0.28 $Y=0.855 $X2=0
+ $Y2=0
cc_136 N_A_27_116#_c_137_n A_269_78# 0.0048076f $X=2.085 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_27_116#_c_137_n A_347_78# 0.0107783f $X=2.085 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_138 N_VPWR_c_197_n N_Y_c_233_n 0.0330222f $X=0.97 $Y=2.035 $X2=0 $Y2=0
cc_139 N_VPWR_c_198_n N_Y_c_233_n 0.0266809f $X=1.97 $Y=2.455 $X2=0 $Y2=0
cc_140 N_VPWR_c_201_n N_Y_c_233_n 0.014552f $X=1.805 $Y=3.33 $X2=0 $Y2=0
cc_141 N_VPWR_c_196_n N_Y_c_233_n 0.0119791f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_142 N_VPWR_M1004_d N_Y_c_243_n 0.0110648f $X=1.77 $Y=1.84 $X2=0 $Y2=0
cc_143 N_VPWR_c_198_n N_Y_c_243_n 0.0232685f $X=1.97 $Y=2.455 $X2=0 $Y2=0
cc_144 N_VPWR_c_198_n Y 0.0282945f $X=1.97 $Y=2.455 $X2=0 $Y2=0
cc_145 N_VPWR_c_203_n Y 0.0217332f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_146 N_VPWR_c_196_n Y 0.0179559f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_147 N_Y_c_231_n N_VGND_c_274_n 0.0221969f $X=2.71 $Y=1.15 $X2=0 $Y2=0
cc_148 N_Y_c_231_n N_VGND_c_275_n 0.0197591f $X=2.71 $Y=1.15 $X2=0 $Y2=0
