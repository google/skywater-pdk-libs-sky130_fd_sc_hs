* File: sky130_fd_sc_hs__ebufn_1.pex.spice
* Created: Tue Sep  1 20:03:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__EBUFN_1%TE_B 1 3 6 10 11 12 14 16 18 19 20 24 25 26
c90 25 0 6.90057e-20 $X=2.03 $Y=2.505
c91 10 0 9.43772e-20 $X=2.68 $Y=1.69
r92 26 36 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.83
r93 26 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.665 $X2=0.59 $Y2=1.665
r94 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.03
+ $Y=2.505 $X2=2.03 $Y2=2.505
r95 19 24 4.82444 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=1.865 $Y=2.505
+ $X2=2.03 $Y2=2.465
r96 19 20 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=1.865 $Y=2.505
+ $X2=0.835 $Y2=2.505
r97 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.75 $Y=2.42
+ $X2=0.835 $Y2=2.505
r98 18 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.75 $Y=2.42 $X2=0.75
+ $Y2=1.83
r99 16 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=2.34
+ $X2=2.03 $Y2=2.505
r100 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.4
r101 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.68 $Y=1.69
+ $X2=2.755 $Y2=1.765
r102 10 11 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.68 $Y=1.69
+ $X2=2.195 $Y2=1.69
r103 8 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=1.765
+ $X2=2.195 $Y2=1.69
r104 8 16 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.12 $Y=1.765
+ $X2=2.12 $Y2=2.34
r105 4 31 38.561 $w=2.98e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.62 $Y=1.5
+ $X2=0.585 $Y2=1.665
r106 4 6 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=0.62 $Y=1.5 $X2=0.62
+ $Y2=0.645
r107 1 31 57.1617 $w=2.98e-07 $l=3.1749e-07 $layer=POLY_cond $X=0.505 $Y=1.945
+ $X2=0.585 $Y2=1.665
r108 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.945
+ $X2=0.505 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_1%A 3 5 7 10 11 15
c36 5 0 9.48915e-20 $X=1.125 $Y=1.945
r37 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.51
+ $Y=1.665 $X2=1.51 $Y2=1.665
r38 11 16 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.51 $Y2=1.665
r39 10 16 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.51
+ $Y2=1.665
r40 9 15 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.215 $Y=1.665
+ $X2=1.51 $Y2=1.665
r41 5 9 68.4907 $w=2.09e-07 $l=2.89828e-07 $layer=POLY_cond $X=1.125 $Y=1.945
+ $X2=1.105 $Y2=1.665
r42 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.125 $Y=1.945
+ $X2=1.125 $Y2=2.44
r43 1 9 41.9691 $w=2.09e-07 $l=1.81659e-07 $layer=POLY_cond $X=1.07 $Y=1.5
+ $X2=1.105 $Y2=1.665
r44 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.07 $Y=1.5 $X2=1.07
+ $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_1%A_27_404# 1 2 7 9 11 14 22 24 25 27 29 33
c61 24 0 9.48915e-20 $X=0.28 $Y=2.165
c62 7 0 9.03051e-20 $X=2.695 $Y=1.295
r63 28 33 35.2787 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.035 $Y=1.24
+ $X2=2.2 $Y2=1.24
r64 27 29 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=1.245
+ $X2=1.87 $Y2=1.245
r65 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.035
+ $Y=1.24 $X2=2.035 $Y2=1.24
r66 24 25 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.165
+ $X2=0.265 $Y2=2
r67 21 22 3.54158 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.53 $Y=1.235
+ $X2=0.307 $Y2=1.235
r68 21 29 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=0.53 $Y=1.235
+ $X2=1.87 $Y2=1.235
r69 16 22 3.0793 $w=3.07e-07 $l=1.74396e-07 $layer=LI1_cond $X=0.17 $Y=1.32
+ $X2=0.307 $Y2=1.235
r70 16 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.17 $Y=1.32
+ $X2=0.17 $Y2=2
r71 12 22 3.0793 $w=3.07e-07 $l=8.5e-08 $layer=LI1_cond $X=0.307 $Y=1.15
+ $X2=0.307 $Y2=1.235
r72 12 14 13.0783 $w=4.43e-07 $l=5.05e-07 $layer=LI1_cond $X=0.307 $Y=1.15
+ $X2=0.307 $Y2=0.645
r73 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.77 $Y=1.185
+ $X2=2.77 $Y2=0.74
r74 7 9 28.2037 $w=2.2e-07 $l=1.42653e-07 $layer=POLY_cond $X=2.695 $Y=1.295
+ $X2=2.77 $Y2=1.185
r75 7 33 144.386 $w=2.2e-07 $l=4.95e-07 $layer=POLY_cond $X=2.695 $Y=1.295
+ $X2=2.2 $Y2=1.295
r76 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.02 $X2=0.28 $Y2=2.165
r77 1 14 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.26
+ $Y=0.37 $X2=0.405 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_1%A_229_74# 1 2 9 11 13 16 18 22 23 24 29 32
+ 35 36 41 42
c92 29 0 9.43772e-20 $X=2.56 $Y=1.32
r93 40 42 12.7871 $w=5.58e-07 $l=5.05e-07 $layer=LI1_cond $X=2.56 $Y=1.6
+ $X2=3.065 $Y2=1.6
r94 40 41 8.50805 $w=5.58e-07 $l=1e-07 $layer=LI1_cond $X=2.56 $Y=1.6 $X2=2.46
+ $Y2=1.6
r95 36 38 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.05 $Y=1.795
+ $X2=2.05 $Y2=2.085
r96 32 42 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.25 $Y=1.485
+ $X2=3.065 $Y2=1.485
r97 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.485 $X2=3.25 $Y2=1.485
r98 29 40 6.84897 $w=2e-07 $l=2.8e-07 $layer=LI1_cond $X=2.56 $Y=1.32 $X2=2.56
+ $Y2=1.6
r99 28 29 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.56 $Y=0.98
+ $X2=2.56 $Y2=1.32
r100 27 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=1.795
+ $X2=2.05 $Y2=1.795
r101 27 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.135 $Y=1.795
+ $X2=2.46 $Y2=1.795
r102 24 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=2.085
+ $X2=2.05 $Y2=2.085
r103 24 35 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.965 $Y=2.085
+ $X2=1.695 $Y2=2.085
r104 22 28 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.46 $Y=0.895
+ $X2=2.56 $Y2=0.98
r105 22 23 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.46 $Y=0.895
+ $X2=1.45 $Y2=0.895
r106 18 35 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.57 $Y=2.125
+ $X2=1.695 $Y2=2.125
r107 18 20 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.57 $Y=2.125
+ $X2=1.355 $Y2=2.125
r108 14 23 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.302 $Y=0.81
+ $X2=1.45 $Y2=0.895
r109 14 16 6.44587 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.302 $Y=0.81
+ $X2=1.302 $Y2=0.645
r110 11 33 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=3.175 $Y=1.765
+ $X2=3.25 $Y2=1.485
r111 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.175 $Y=1.765
+ $X2=3.175 $Y2=2.4
r112 7 33 38.6072 $w=2.91e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.16 $Y=1.32
+ $X2=3.25 $Y2=1.485
r113 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.16 $Y=1.32 $X2=3.16
+ $Y2=0.74
r114 2 20 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.02 $X2=1.355 $Y2=2.165
r115 1 16 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.37 $X2=1.285 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_1%VPWR 1 2 11 15 19 21 31 32 35 38
c46 32 0 6.90057e-20 $X=3.6 $Y=3.33
c47 15 0 9.03051e-20 $X=2.53 $Y=2.135
r48 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 32 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.53 $Y2=3.33
r53 29 31 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 25 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r58 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 22 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r60 22 24 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 21 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.53 $Y2=3.33
r62 21 27 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 19 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r64 19 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.53 $Y=2.135
+ $X2=2.53 $Y2=2.815
r66 13 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=3.33
r67 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=2.815
r68 9 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r69 9 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.925
r70 2 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.84 $X2=2.53 $Y2=2.815
r71 2 15 400 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.84 $X2=2.53 $Y2=2.135
r72 1 11 600 $w=1.7e-07 $l=1.01573e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.02 $X2=0.815 $Y2=2.925
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_1%Z 1 2 9 14 15 16 17 21
r25 17 27 10.6778 $w=5.43e-07 $l=2.05e-07 $layer=LI1_cond $X=3.482 $Y=0.925
+ $X2=3.482 $Y2=1.13
r26 16 17 8.12016 $w=5.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.482 $Y=0.555
+ $X2=3.482 $Y2=0.925
r27 16 21 0.877856 $w=5.43e-07 $l=4e-08 $layer=LI1_cond $X=3.482 $Y=0.555
+ $X2=3.482 $Y2=0.515
r28 15 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.82 $X2=3.67
+ $Y2=1.13
r29 14 15 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=1.985
+ $X2=3.495 $Y2=1.82
r30 7 14 2.18514 $w=5.18e-07 $l=9.5e-08 $layer=LI1_cond $X=3.495 $Y=2.08
+ $X2=3.495 $Y2=1.985
r31 7 9 16.9061 $w=5.18e-07 $l=7.35e-07 $layer=LI1_cond $X=3.495 $Y=2.08
+ $X2=3.495 $Y2=2.815
r32 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.25
+ $Y=1.84 $X2=3.4 $Y2=1.985
r33 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.25
+ $Y=1.84 $X2=3.4 $Y2=2.815
r34 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.235
+ $Y=0.37 $X2=3.375 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__EBUFN_1%VGND 1 2 11 15 17 19 29 30 33 36
r32 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r33 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r34 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r35 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r36 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.555
+ $Y2=0
r37 27 29 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=3.6
+ $Y2=0
r38 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r39 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r41 22 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r42 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 20 33 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.842
+ $Y2=0
r44 20 22 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.2
+ $Y2=0
r45 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.555
+ $Y2=0
r46 19 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.16
+ $Y2=0
r47 17 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r48 17 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r49 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=0.085
+ $X2=2.555 $Y2=0
r50 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.555 $Y=0.085
+ $X2=2.555 $Y2=0.535
r51 9 33 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0
r52 9 11 22.6445 $w=2.83e-07 $l=5.6e-07 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0.645
r53 2 15 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=2.41
+ $Y=0.37 $X2=2.555 $Y2=0.535
r54 1 11 182 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_NDIFF $count=1 $X=0.695
+ $Y=0.37 $X2=0.845 $Y2=0.645
.ends

