# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__o221ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o221ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.300000 3.715000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.350000 2.775000 1.680000 ;
        RECT 2.525000 1.680000 2.775000 2.890000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.350000 1.635000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.875000 1.350000 2.275000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.011700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.445000 0.960000 ;
        RECT 0.115000 0.960000 0.775000 1.130000 ;
        RECT 0.325000 1.950000 2.355000 2.120000 ;
        RECT 0.325000 2.120000 0.575000 2.980000 ;
        RECT 0.605000 1.130000 0.775000 1.950000 ;
        RECT 2.025000 2.120000 2.355000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.840000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 4.030000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.615000  0.350000 2.005000 0.520000 ;
      RECT 0.615000  0.520000 0.945000 0.770000 ;
      RECT 0.745000  2.290000 1.560000 3.245000 ;
      RECT 1.175000  0.800000 1.505000 1.010000 ;
      RECT 1.175000  1.010000 3.725000 1.130000 ;
      RECT 1.175000  1.130000 2.505000 1.180000 ;
      RECT 1.675000  0.520000 2.005000 0.795000 ;
      RECT 2.175000  0.350000 2.505000 0.960000 ;
      RECT 2.175000  0.960000 3.725000 1.010000 ;
      RECT 2.675000  0.085000 3.225000 0.790000 ;
      RECT 3.165000  1.950000 3.495000 3.245000 ;
      RECT 3.395000  0.350000 3.725000 0.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o221ai_1
END LIBRARY
