* File: sky130_fd_sc_hs__dlrtp_1.spice
* Created: Tue Sep  1 20:02:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlrtp_1.pex.spice"
.subckt sky130_fd_sc_hs__dlrtp_1  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_D_M1017_g N_A_27_424#_M1017_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.125093 AS=0.15675 PD=1.00194 PS=1.67 NRD=34.356 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1002 N_A_216_424#_M1002_d N_GATE_M1002_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.168307 PD=2.05 PS=1.34806 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_216_424#_M1010_g N_A_363_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.136954 AS=0.32225 PD=1.17971 PS=2.64 NRD=4.86 NRS=61.692 M=1
+ R=4.93333 SA=75000.3 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1018 A_565_74# N_A_27_424#_M1018_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.118446 PD=0.88 PS=1.02029 NRD=12.18 NRS=9.372 M=1 R=4.26667
+ SA=75000.8 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1019 N_A_643_74#_M1019_d N_A_363_74#_M1019_g A_565_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.175517 AS=0.0768 PD=1.35245 PS=0.88 NRD=11.244 NRS=12.18 M=1
+ R=4.26667 SA=75001.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1006 A_769_74# N_A_216_424#_M1006_g N_A_643_74#_M1019_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.115183 PD=0.66 PS=0.887547 NRD=18.564 NRS=41.424 M=1
+ R=2.8 SA=75001.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_817_48#_M1007_g A_769_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_1045_74# N_A_643_74#_M1015_g N_A_817_48#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_RESET_B_M1003_g A_1045_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.0888 PD=1.1 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_Q_M1013_d N_A_817_48#_M1013_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1332 PD=2.05 PS=1.1 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_A_27_424#_M1012_s VPB PSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.2478 PD=1.19 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1009 N_A_216_424#_M1009_d N_GATE_M1009_g N_VPWR_M1012_d VPB PSHORT L=0.15
+ W=0.84 AD=0.43935 AS=0.147 PD=2.87 PS=1.19 NRD=32.8202 NRS=2.3443 M=1 R=5.6
+ SA=75000.7 SB=75000.4 A=0.126 P=1.98 MULT=1
MM1011 N_VPWR_M1011_d N_A_216_424#_M1011_g N_A_363_74#_M1011_s VPB PSHORT L=0.15
+ W=0.84 AD=0.18973 AS=0.2478 PD=1.30565 PS=2.27 NRD=28.1316 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1000 A_568_392# N_A_27_424#_M1000_g N_VPWR_M1011_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.22587 PD=1.27 PS=1.55435 NRD=15.7403 NRS=6.8753 M=1 R=6.66667
+ SA=75000.7 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1008 N_A_643_74#_M1008_d N_A_216_424#_M1008_g A_568_392# VPB PSHORT L=0.15 W=1
+ AD=0.234366 AS=0.135 PD=1.9507 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.1 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1005 A_759_508# N_A_363_74#_M1005_g N_A_643_74#_M1008_d VPB PSHORT L=0.15
+ W=0.42 AD=0.10605 AS=0.0984338 PD=0.925 PS=0.819296 NRD=92.6294 NRS=46.886 M=1
+ R=2.8 SA=75001.6 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_817_48#_M1001_g A_759_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.121238 AS=0.10605 PD=0.952394 PS=0.925 NRD=77.3816 NRS=92.6294 M=1 R=2.8
+ SA=75002.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1016 N_A_817_48#_M1016_d N_A_643_74#_M1016_g N_VPWR_M1001_d VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.288662 PD=1.35 PS=2.26761 NRD=11.8003 NRS=32.4853 M=1
+ R=6.66667 SA=75001.4 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_RESET_B_M1014_g N_A_817_48#_M1016_d VPB PSHORT L=0.15
+ W=1 AD=0.21783 AS=0.175 PD=1.46226 PS=1.35 NRD=11.8003 NRS=1.9503 M=1
+ R=6.66667 SA=75001.9 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1004 N_Q_M1004_d N_A_817_48#_M1004_g N_VPWR_M1014_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.24397 PD=2.83 PS=1.63774 NRD=1.7533 NRS=15.8191 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.9966 P=18.16
c_860 A_568_392# 0 1.90301e-19 $X=2.84 $Y=1.96
c_961 A_565_74# 0 5.47968e-20 $X=2.825 $Y=0.37
*
.include "sky130_fd_sc_hs__dlrtp_1.pxi.spice"
*
.ends
*
*
