* File: sky130_fd_sc_hs__einvn_2.spice
* Created: Thu Aug 27 20:44:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__einvn_2.pex.spice"
.subckt sky130_fd_sc_hs__einvn_2  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1009 N_A_115_464#_M1009_d N_TE_B_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_115_464#_M1000_g N_A_231_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1000_d N_A_115_464#_M1003_g N_A_231_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_231_74#_M1003_s N_A_M1001_g N_Z_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.10545 PD=1.02 PS=1.025 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_A_231_74#_M1008_d N_A_M1008_g N_Z_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1995 AS=0.10545 PD=2.08 PS=1.025 NRD=0 NRS=0.804 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_115_464#_M1007_d N_TE_B_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15
+ W=0.64 AD=0.1856 AS=0.1856 PD=1.86 PS=1.86 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_TE_B_M1002_g N_A_227_368#_M1002_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1002_d N_TE_B_M1004_g N_A_227_368#_M1004_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1005 N_Z_M1005_d N_A_M1005_g N_A_227_368#_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_Z_M1005_d N_A_M1006_g N_A_227_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__einvn_2.pxi.spice"
*
.ends
*
*
