* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__and3_4 A B C VGND VNB VPB VPWR X
X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 VPWR B a_83_260# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 a_83_260# C VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X4 VGND C a_489_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_686_74# B a_489_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 a_83_260# A a_686_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_489_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_489_74# B a_686_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_83_260# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VPWR C a_83_260# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X18 a_686_74# A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
