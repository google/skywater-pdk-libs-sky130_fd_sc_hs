# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a32oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a32oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.180000 2.775000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.375000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.785000 1.180000 6.115000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.180000 2.275000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 1.090000 1.630000 ;
        RECT 0.125000 1.630000 0.355000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.192800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.800000 3.235000 1.890000 ;
        RECT 0.615000 1.890000 1.945000 1.970000 ;
        RECT 0.615000 1.970000 0.945000 2.735000 ;
        RECT 1.455000 0.595000 1.785000 0.840000 ;
        RECT 1.455000 0.840000 3.205000 1.010000 ;
        RECT 1.615000 1.720000 3.235000 1.800000 ;
        RECT 1.615000 1.970000 1.945000 2.735000 ;
        RECT 3.005000 1.010000 3.205000 1.235000 ;
        RECT 3.005000 1.235000 3.235000 1.720000 ;
        RECT 3.015000 0.595000 3.205000 0.840000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.960000 ;
      RECT 0.115000  0.960000 1.275000 1.130000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.400000 3.075000 ;
      RECT 0.545000  0.085000 0.875000 0.790000 ;
      RECT 1.105000  0.255000 2.285000 0.425000 ;
      RECT 1.105000  0.425000 1.275000 0.960000 ;
      RECT 1.115000  2.140000 1.445000 2.905000 ;
      RECT 1.955000  0.425000 2.285000 0.670000 ;
      RECT 2.115000  2.060000 4.875000 2.120000 ;
      RECT 2.115000  2.120000 3.735000 2.230000 ;
      RECT 2.115000  2.230000 2.400000 2.905000 ;
      RECT 2.515000  0.255000 4.705000 0.425000 ;
      RECT 2.515000  0.425000 2.845000 0.670000 ;
      RECT 2.570000  2.400000 3.280000 3.245000 ;
      RECT 3.375000  0.425000 3.705000 1.130000 ;
      RECT 3.405000  1.950000 4.875000 2.060000 ;
      RECT 3.450000  2.230000 3.735000 2.980000 ;
      RECT 3.875000  0.595000 4.205000 1.010000 ;
      RECT 3.875000  1.010000 5.615000 1.180000 ;
      RECT 3.905000  2.290000 4.250000 3.245000 ;
      RECT 4.375000  0.425000 4.705000 0.840000 ;
      RECT 4.420000  2.120000 4.875000 2.980000 ;
      RECT 4.545000  1.720000 5.875000 1.890000 ;
      RECT 4.545000  1.890000 4.875000 1.950000 ;
      RECT 4.935000  0.085000 5.185000 0.840000 ;
      RECT 5.045000  2.060000 5.375000 3.245000 ;
      RECT 5.365000  0.350000 5.615000 1.010000 ;
      RECT 5.545000  1.890000 5.875000 2.980000 ;
      RECT 5.795000  0.085000 6.125000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__a32oi_2
END LIBRARY
