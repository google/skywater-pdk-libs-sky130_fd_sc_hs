* File: sky130_fd_sc_hs__a21o_4.spice
* Created: Tue Sep  1 19:49:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a21o_4.pex.spice"
.subckt sky130_fd_sc_hs__a21o_4  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_X_M1006_d N_A_91_48#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1006_d N_A_91_48#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1012_d N_A_91_48#_M1012_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1012_d N_A_91_48#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.130894 PD=1.02 PS=1.15826 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1011 N_A_91_48#_M1011_d N_B1_M1011_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.113206 PD=0.92 PS=1.00174 NRD=0 NRS=11.244 M=1 R=4.26667
+ SA=75002 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1017 N_A_91_48#_M1011_d N_B1_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_700_74#_M1009_d N_A1_M1009_g N_A_91_48#_M1009_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1015 N_A_700_74#_M1015_d N_A1_M1015_g N_A_91_48#_M1009_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_700_74#_M1015_d N_A2_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1014 N_A_700_74#_M1014_d N_A2_M1014_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_X_M1002_d N_A_91_48#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1004 N_X_M1002_d N_A_91_48#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1018 N_X_M1018_d N_A_91_48#_M1018_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1019 N_X_M1018_d N_A_91_48#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_503_392#_M1000_d N_B1_M1000_g N_A_91_48#_M1000_s VPB PSHORT L=0.15
+ W=1 AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1016 N_A_503_392#_M1016_d N_B1_M1016_g N_A_91_48#_M1000_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75002 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_503_392#_M1016_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1003_d N_A1_M1005_g N_A_503_392#_M1005_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_503_392#_M1005_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1007_d N_A2_M1008_g N_A_503_392#_M1008_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_hs__a21o_4.pxi.spice"
*
.ends
*
*
