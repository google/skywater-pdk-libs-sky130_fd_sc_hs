* File: sky130_fd_sc_hs__o21ba_4.pxi.spice
* Created: Thu Aug 27 20:58:38 2020
* 
x_PM_SKY130_FD_SC_HS__O21BA_4%B1_N N_B1_N_c_115_n N_B1_N_M1016_g N_B1_N_c_116_n
+ N_B1_N_M1021_g B1_N PM_SKY130_FD_SC_HS__O21BA_4%B1_N
x_PM_SKY130_FD_SC_HS__O21BA_4%A_193_48# N_A_193_48#_M1007_d N_A_193_48#_M1000_d
+ N_A_193_48#_M1008_d N_A_193_48#_M1002_g N_A_193_48#_c_160_n
+ N_A_193_48#_M1011_g N_A_193_48#_M1005_g N_A_193_48#_c_161_n
+ N_A_193_48#_M1012_g N_A_193_48#_M1013_g N_A_193_48#_c_162_n
+ N_A_193_48#_M1014_g N_A_193_48#_M1020_g N_A_193_48#_c_163_n
+ N_A_193_48#_M1017_g N_A_193_48#_c_152_n N_A_193_48#_c_153_n
+ N_A_193_48#_c_154_n N_A_193_48#_c_155_n N_A_193_48#_c_156_n
+ N_A_193_48#_c_177_p N_A_193_48#_c_157_n N_A_193_48#_c_164_n
+ N_A_193_48#_c_165_n N_A_193_48#_c_207_p N_A_193_48#_c_158_n
+ N_A_193_48#_c_166_n N_A_193_48#_c_159_n PM_SKY130_FD_SC_HS__O21BA_4%A_193_48#
x_PM_SKY130_FD_SC_HS__O21BA_4%A_27_368# N_A_27_368#_M1021_s N_A_27_368#_M1016_s
+ N_A_27_368#_c_318_n N_A_27_368#_M1000_g N_A_27_368#_M1007_g
+ N_A_27_368#_c_319_n N_A_27_368#_M1001_g N_A_27_368#_M1019_g
+ N_A_27_368#_c_313_n N_A_27_368#_c_320_n N_A_27_368#_c_321_n
+ N_A_27_368#_c_331_n N_A_27_368#_c_322_n N_A_27_368#_c_314_n
+ N_A_27_368#_c_323_n N_A_27_368#_c_315_n N_A_27_368#_c_325_n
+ N_A_27_368#_c_316_n N_A_27_368#_c_317_n PM_SKY130_FD_SC_HS__O21BA_4%A_27_368#
x_PM_SKY130_FD_SC_HS__O21BA_4%A2 N_A2_c_414_n N_A2_M1008_g N_A2_M1003_g
+ N_A2_c_415_n N_A2_M1015_g N_A2_M1009_g A2 A2 A2 N_A2_c_413_n
+ PM_SKY130_FD_SC_HS__O21BA_4%A2
x_PM_SKY130_FD_SC_HS__O21BA_4%A1 N_A1_M1006_g N_A1_c_470_n N_A1_M1004_g
+ N_A1_c_471_n N_A1_c_472_n N_A1_c_473_n N_A1_c_474_n N_A1_c_479_n N_A1_M1018_g
+ N_A1_M1010_g A1 PM_SKY130_FD_SC_HS__O21BA_4%A1
x_PM_SKY130_FD_SC_HS__O21BA_4%VPWR N_VPWR_M1016_d N_VPWR_M1012_s N_VPWR_M1017_s
+ N_VPWR_M1001_s N_VPWR_M1018_s N_VPWR_c_540_n N_VPWR_c_541_n N_VPWR_c_542_n
+ N_VPWR_c_543_n N_VPWR_c_544_n VPWR N_VPWR_c_545_n N_VPWR_c_546_n
+ N_VPWR_c_547_n N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n
+ N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_539_n PM_SKY130_FD_SC_HS__O21BA_4%VPWR
x_PM_SKY130_FD_SC_HS__O21BA_4%X N_X_M1002_s N_X_M1013_s N_X_M1011_d N_X_M1014_d
+ N_X_c_617_n N_X_c_623_n N_X_c_618_n N_X_c_619_n N_X_c_620_n X X N_X_c_626_n X
+ N_X_c_622_n PM_SKY130_FD_SC_HS__O21BA_4%X
x_PM_SKY130_FD_SC_HS__O21BA_4%A_892_392# N_A_892_392#_M1004_d
+ N_A_892_392#_M1015_s N_A_892_392#_c_673_n N_A_892_392#_c_669_n
+ N_A_892_392#_c_670_n N_A_892_392#_c_671_n
+ PM_SKY130_FD_SC_HS__O21BA_4%A_892_392#
x_PM_SKY130_FD_SC_HS__O21BA_4%VGND N_VGND_M1021_d N_VGND_M1005_d N_VGND_M1020_d
+ N_VGND_M1006_s N_VGND_M1009_d N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n
+ N_VGND_c_703_n N_VGND_c_704_n N_VGND_c_705_n N_VGND_c_706_n VGND
+ N_VGND_c_707_n N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n
+ N_VGND_c_712_n N_VGND_c_713_n N_VGND_c_714_n N_VGND_c_715_n
+ PM_SKY130_FD_SC_HS__O21BA_4%VGND
x_PM_SKY130_FD_SC_HS__O21BA_4%A_618_94# N_A_618_94#_M1007_s N_A_618_94#_M1019_s
+ N_A_618_94#_M1003_s N_A_618_94#_M1010_d N_A_618_94#_c_800_n
+ N_A_618_94#_c_791_n N_A_618_94#_c_792_n N_A_618_94#_c_793_n
+ N_A_618_94#_c_794_n N_A_618_94#_c_795_n N_A_618_94#_c_796_n
+ N_A_618_94#_c_797_n N_A_618_94#_c_798_n N_A_618_94#_c_799_n
+ PM_SKY130_FD_SC_HS__O21BA_4%A_618_94#
cc_1 VNB N_B1_N_c_115_n 0.0438568f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_B1_N_c_116_n 0.0222506f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.22
cc_3 VNB B1_N 0.00980764f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_193_48#_M1002_g 0.0210367f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.365
cc_5 VNB N_A_193_48#_M1005_g 0.0199949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_193_48#_M1013_g 0.020485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_193_48#_M1020_g 0.0235858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_193_48#_c_152_n 0.0209991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_193_48#_c_153_n 0.0190649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_193_48#_c_154_n 0.0166372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_193_48#_c_155_n 0.0034847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_193_48#_c_156_n 0.0206699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_193_48#_c_157_n 0.00158703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_193_48#_c_158_n 0.0112053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_193_48#_c_159_n 0.109811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_368#_M1007_g 0.0421943f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.365
cc_17 VNB N_A_27_368#_M1019_g 0.0367602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_368#_c_313_n 0.0222049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_368#_c_314_n 0.0079873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_368#_c_315_n 0.0300846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_368#_c_316_n 5.55182e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_368#_c_317_n 0.0117632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_M1003_g 0.0196921f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.74
cc_24 VNB N_A2_M1009_g 0.0180242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB A2 0.0144679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_413_n 0.0248587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_M1006_g 0.0327623f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.22
cc_28 VNB N_A1_c_470_n 0.0163721f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.74
cc_29 VNB N_A1_c_471_n 0.0975279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_c_472_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.385
cc_31 VNB N_A1_c_473_n 0.00843327f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_32 VNB N_A1_c_474_n 0.0143086f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_33 VNB N_A1_M1010_g 0.0360452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB A1 0.00447618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_539_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_617_n 0.00202189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_618_n 0.00629496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_619_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_620_n 0.00111459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB X 7.86953e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_622_n 0.00286244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_700_n 0.00587905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_701_n 0.00412957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_702_n 0.00722278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_703_n 0.0100107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_704_n 0.00760342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_705_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_706_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_707_n 0.0157739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_708_n 0.0469424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_709_n 0.0160823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_710_n 0.0195709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_711_n 0.350143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_712_n 0.0258092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_713_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_714_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_715_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_618_94#_c_791_n 0.00431549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_618_94#_c_792_n 0.00135951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_618_94#_c_793_n 0.00127304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_618_94#_c_794_n 0.00363185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_618_94#_c_795_n 0.0020675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_618_94#_c_796_n 0.0130457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_618_94#_c_797_n 0.0231872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_618_94#_c_798_n 0.00541364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_618_94#_c_799_n 0.00177818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VPB N_B1_N_c_115_n 0.0291938f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_68 VPB N_A_193_48#_c_160_n 0.0155966f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_69 VPB N_A_193_48#_c_161_n 0.0148723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_193_48#_c_162_n 0.0148883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_193_48#_c_163_n 0.0178512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_193_48#_c_164_n 0.00977712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_193_48#_c_165_n 0.00110611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_193_48#_c_166_n 0.00347163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_193_48#_c_159_n 0.0272311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_27_368#_c_318_n 0.0169557f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_77 VPB N_A_27_368#_c_319_n 0.0160349f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_78 VPB N_A_27_368#_c_320_n 0.0153183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_27_368#_c_321_n 0.0195781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_27_368#_c_322_n 0.0023962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_27_368#_c_323_n 0.01385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_27_368#_c_315_n 0.00777552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_27_368#_c_325_n 0.00723806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_27_368#_c_316_n 0.00482872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_27_368#_c_317_n 0.0625278f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A2_c_414_n 0.0147804f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_87 VPB N_A2_c_415_n 0.0148371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB A2 0.0119519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A2_c_413_n 0.03352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A1_c_470_n 0.0340202f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.74
cc_91 VPB N_A1_c_474_n 0.00848991f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.385
cc_92 VPB N_A1_c_479_n 0.0266121f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.365
cc_93 VPB A1 0.00323349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_540_n 0.00639038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_541_n 0.00261656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_542_n 0.00936969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_543_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_544_n 0.051587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_545_n 0.0189171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_546_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_547_n 0.0215473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_548_n 0.0387727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_549_n 0.00710329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_550_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_551_n 0.017758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_552_n 0.024435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_553_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_539_n 0.073215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_X_c_623_n 0.00516914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB X 0.00146868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_892_392#_c_669_n 0.00431993f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.385
cc_112 VPB N_A_892_392#_c_670_n 0.00217954f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.365
cc_113 VPB N_A_892_392#_c_671_n 0.00268696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 N_B1_N_c_115_n N_A_193_48#_M1002_g 0.0212371f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_B1_N_c_116_n N_A_193_48#_M1002_g 0.0168899f $X=0.525 $Y=1.22 $X2=0
+ $Y2=0
cc_116 B1_N N_A_193_48#_M1002_g 0.00324428f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B1_N_c_115_n N_A_193_48#_c_160_n 0.0318301f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_B1_N_c_115_n N_A_193_48#_c_159_n 0.00756852f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_B1_N_c_116_n N_A_27_368#_c_313_n 0.00581235f $X=0.525 $Y=1.22 $X2=0
+ $Y2=0
cc_120 N_B1_N_c_115_n N_A_27_368#_c_320_n 0.0080039f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_121 N_B1_N_c_115_n N_A_27_368#_c_321_n 0.00675288f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_B1_N_c_115_n N_A_27_368#_c_331_n 0.0134961f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_B1_N_c_116_n N_A_27_368#_c_314_n 0.00232983f $X=0.525 $Y=1.22 $X2=0
+ $Y2=0
cc_124 B1_N N_A_27_368#_c_314_n 0.00294872f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_125 N_B1_N_c_115_n N_A_27_368#_c_323_n 0.00478733f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_126 B1_N N_A_27_368#_c_323_n 0.00107809f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_N_c_115_n N_A_27_368#_c_315_n 0.0152937f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_B1_N_c_116_n N_A_27_368#_c_315_n 0.00346495f $X=0.525 $Y=1.22 $X2=0
+ $Y2=0
cc_129 B1_N N_A_27_368#_c_315_n 0.0284252f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_130 N_B1_N_c_115_n N_A_27_368#_c_325_n 2.24111e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_B1_N_c_115_n N_VPWR_c_540_n 0.00483983f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_132 N_B1_N_c_115_n N_VPWR_c_545_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_133 N_B1_N_c_115_n N_VPWR_c_539_n 0.00440701f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_134 N_B1_N_c_115_n X 0.0012955f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_135 N_B1_N_c_115_n N_X_c_626_n 0.00128628f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_136 N_B1_N_c_115_n N_X_c_622_n 2.26341e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_137 B1_N N_X_c_622_n 0.0185939f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_138 N_B1_N_c_115_n N_VGND_c_700_n 7.44677e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_139 N_B1_N_c_116_n N_VGND_c_700_n 0.00674192f $X=0.525 $Y=1.22 $X2=0 $Y2=0
cc_140 B1_N N_VGND_c_700_n 0.0160286f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_141 N_B1_N_c_116_n N_VGND_c_711_n 0.0082465f $X=0.525 $Y=1.22 $X2=0 $Y2=0
cc_142 N_B1_N_c_116_n N_VGND_c_712_n 0.00434272f $X=0.525 $Y=1.22 $X2=0 $Y2=0
cc_143 N_A_193_48#_c_166_n N_A_27_368#_c_318_n 0.00689099f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_144 N_A_193_48#_c_153_n N_A_27_368#_M1007_g 0.00845542f $X=2.895 $Y=1.29
+ $X2=0 $Y2=0
cc_145 N_A_193_48#_c_154_n N_A_27_368#_M1007_g 0.00964849f $X=3.5 $Y=0.34 $X2=0
+ $Y2=0
cc_146 N_A_193_48#_c_156_n N_A_27_368#_M1007_g 0.0129483f $X=3.66 $Y=1.375 $X2=0
+ $Y2=0
cc_147 N_A_193_48#_c_177_p N_A_27_368#_M1007_g 0.00612159f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_148 N_A_193_48#_c_157_n N_A_27_368#_M1007_g 0.00364839f $X=3.745 $Y=1.95
+ $X2=0 $Y2=0
cc_149 N_A_193_48#_c_158_n N_A_27_368#_M1007_g 0.00518238f $X=2.895 $Y=1.455
+ $X2=0 $Y2=0
cc_150 N_A_193_48#_c_164_n N_A_27_368#_c_319_n 0.00725299f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_151 N_A_193_48#_c_166_n N_A_27_368#_c_319_n 0.0177723f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_152 N_A_193_48#_c_154_n N_A_27_368#_M1019_g 0.00312284f $X=3.5 $Y=0.34 $X2=0
+ $Y2=0
cc_153 N_A_193_48#_c_156_n N_A_27_368#_M1019_g 0.00586411f $X=3.66 $Y=1.375
+ $X2=0 $Y2=0
cc_154 N_A_193_48#_c_177_p N_A_27_368#_M1019_g 0.00621111f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_155 N_A_193_48#_c_157_n N_A_27_368#_M1019_g 0.00355214f $X=3.745 $Y=1.95
+ $X2=0 $Y2=0
cc_156 N_A_193_48#_c_160_n N_A_27_368#_c_321_n 5.6504e-19 $X=1.055 $Y=1.765
+ $X2=0 $Y2=0
cc_157 N_A_193_48#_c_160_n N_A_27_368#_c_331_n 0.0154267f $X=1.055 $Y=1.765
+ $X2=0 $Y2=0
cc_158 N_A_193_48#_c_161_n N_A_27_368#_c_331_n 0.0117914f $X=1.505 $Y=1.765
+ $X2=0 $Y2=0
cc_159 N_A_193_48#_c_162_n N_A_27_368#_c_331_n 0.0117914f $X=1.955 $Y=1.765
+ $X2=0 $Y2=0
cc_160 N_A_193_48#_c_163_n N_A_27_368#_c_331_n 0.0178278f $X=2.405 $Y=1.765
+ $X2=0 $Y2=0
cc_161 N_A_193_48#_c_166_n N_A_27_368#_c_331_n 0.0137304f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_162 N_A_193_48#_c_163_n N_A_27_368#_c_322_n 0.00878392f $X=2.405 $Y=1.765
+ $X2=0 $Y2=0
cc_163 N_A_193_48#_c_166_n N_A_27_368#_c_322_n 0.0280237f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_164 N_A_193_48#_c_160_n N_A_27_368#_c_323_n 0.00198831f $X=1.055 $Y=1.765
+ $X2=0 $Y2=0
cc_165 N_A_193_48#_c_163_n N_A_27_368#_c_316_n 0.00295122f $X=2.405 $Y=1.765
+ $X2=0 $Y2=0
cc_166 N_A_193_48#_c_156_n N_A_27_368#_c_316_n 0.025164f $X=3.66 $Y=1.375 $X2=0
+ $Y2=0
cc_167 N_A_193_48#_c_157_n N_A_27_368#_c_316_n 0.0229207f $X=3.745 $Y=1.95 $X2=0
+ $Y2=0
cc_168 N_A_193_48#_c_166_n N_A_27_368#_c_316_n 7.23724e-19 $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_169 N_A_193_48#_c_159_n N_A_27_368#_c_316_n 0.0020839f $X=2.34 $Y=1.527 $X2=0
+ $Y2=0
cc_170 N_A_193_48#_c_163_n N_A_27_368#_c_317_n 0.00230301f $X=2.405 $Y=1.765
+ $X2=0 $Y2=0
cc_171 N_A_193_48#_c_156_n N_A_27_368#_c_317_n 0.00645374f $X=3.66 $Y=1.375
+ $X2=0 $Y2=0
cc_172 N_A_193_48#_c_157_n N_A_27_368#_c_317_n 0.0148458f $X=3.745 $Y=1.95 $X2=0
+ $Y2=0
cc_173 N_A_193_48#_c_164_n N_A_27_368#_c_317_n 0.00804416f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_174 N_A_193_48#_c_166_n N_A_27_368#_c_317_n 0.00954859f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_175 N_A_193_48#_c_159_n N_A_27_368#_c_317_n 0.00168876f $X=2.34 $Y=1.527
+ $X2=0 $Y2=0
cc_176 N_A_193_48#_c_164_n N_A2_c_414_n 0.016535f $X=4.975 $Y=2.125 $X2=-0.19
+ $Y2=-0.245
cc_177 N_A_193_48#_c_207_p N_A2_c_414_n 0.00440627f $X=5.06 $Y=2.57 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A_193_48#_c_165_n N_A2_c_415_n 0.00157886f $X=5.06 $Y=2.3 $X2=0 $Y2=0
cc_179 N_A_193_48#_c_207_p N_A2_c_415_n 0.00165372f $X=5.06 $Y=2.57 $X2=0 $Y2=0
cc_180 N_A_193_48#_c_164_n A2 0.0100261f $X=4.975 $Y=2.125 $X2=0 $Y2=0
cc_181 N_A_193_48#_c_165_n A2 0.0143367f $X=5.06 $Y=2.3 $X2=0 $Y2=0
cc_182 N_A_193_48#_c_164_n N_A2_c_413_n 0.00230545f $X=4.975 $Y=2.125 $X2=0
+ $Y2=0
cc_183 N_A_193_48#_c_165_n N_A2_c_413_n 0.00423635f $X=5.06 $Y=2.3 $X2=0 $Y2=0
cc_184 N_A_193_48#_c_154_n N_A1_M1006_g 0.00179591f $X=3.5 $Y=0.34 $X2=0 $Y2=0
cc_185 N_A_193_48#_c_156_n N_A1_M1006_g 7.47639e-19 $X=3.66 $Y=1.375 $X2=0 $Y2=0
cc_186 N_A_193_48#_c_177_p N_A1_M1006_g 6.35849e-19 $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_187 N_A_193_48#_c_157_n N_A1_c_470_n 0.00122424f $X=3.745 $Y=1.95 $X2=0 $Y2=0
cc_188 N_A_193_48#_c_164_n N_A1_c_470_n 0.0278886f $X=4.975 $Y=2.125 $X2=0 $Y2=0
cc_189 N_A_193_48#_c_166_n N_A1_c_470_n 8.72368e-19 $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_190 N_A_193_48#_c_156_n A1 4.2002e-19 $X=3.66 $Y=1.375 $X2=0 $Y2=0
cc_191 N_A_193_48#_c_157_n A1 0.013357f $X=3.745 $Y=1.95 $X2=0 $Y2=0
cc_192 N_A_193_48#_c_164_n A1 0.0398385f $X=4.975 $Y=2.125 $X2=0 $Y2=0
cc_193 N_A_193_48#_c_164_n N_VPWR_M1001_s 0.00510692f $X=4.975 $Y=2.125 $X2=0
+ $Y2=0
cc_194 N_A_193_48#_c_160_n N_VPWR_c_540_n 0.00855671f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_193_48#_c_161_n N_VPWR_c_540_n 0.0010638f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_193_48#_c_160_n N_VPWR_c_541_n 0.00106466f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_193_48#_c_161_n N_VPWR_c_541_n 0.00840438f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_193_48#_c_162_n N_VPWR_c_541_n 0.00838241f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A_193_48#_c_163_n N_VPWR_c_541_n 0.00106604f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_193_48#_c_164_n N_VPWR_c_542_n 0.0262543f $X=4.975 $Y=2.125 $X2=0
+ $Y2=0
cc_201 N_A_193_48#_c_166_n N_VPWR_c_542_n 0.0336225f $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_202 N_A_193_48#_c_160_n N_VPWR_c_546_n 0.00413917f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_193_48#_c_161_n N_VPWR_c_546_n 0.00413917f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A_193_48#_c_166_n N_VPWR_c_547_n 0.0110241f $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_205 N_A_193_48#_c_162_n N_VPWR_c_551_n 0.00413917f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_193_48#_c_163_n N_VPWR_c_551_n 0.00413917f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_193_48#_c_162_n N_VPWR_c_552_n 0.00105871f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_193_48#_c_163_n N_VPWR_c_552_n 0.00991572f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_193_48#_c_166_n N_VPWR_c_552_n 0.0142559f $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_210 N_A_193_48#_c_160_n N_VPWR_c_539_n 0.00398641f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_A_193_48#_c_161_n N_VPWR_c_539_n 0.00398641f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_A_193_48#_c_162_n N_VPWR_c_539_n 0.00398641f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A_193_48#_c_163_n N_VPWR_c_539_n 0.00397108f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A_193_48#_c_166_n N_VPWR_c_539_n 0.00909194f $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_215 N_A_193_48#_M1002_g N_X_c_617_n 3.77529e-19 $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_193_48#_M1005_g N_X_c_617_n 0.00305913f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_193_48#_c_161_n N_X_c_623_n 0.017138f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_193_48#_c_162_n N_X_c_623_n 0.0153034f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_193_48#_c_163_n N_X_c_623_n 0.0190908f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_193_48#_c_152_n N_X_c_623_n 0.0600869f $X=2.81 $Y=1.455 $X2=0 $Y2=0
cc_221 N_A_193_48#_c_159_n N_X_c_623_n 0.0201796f $X=2.34 $Y=1.527 $X2=0 $Y2=0
cc_222 N_A_193_48#_M1005_g N_X_c_618_n 0.0147036f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_193_48#_M1013_g N_X_c_618_n 0.0119326f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_193_48#_c_152_n N_X_c_618_n 0.0559114f $X=2.81 $Y=1.455 $X2=0 $Y2=0
cc_225 N_A_193_48#_c_159_n N_X_c_618_n 0.00457162f $X=2.34 $Y=1.527 $X2=0 $Y2=0
cc_226 N_A_193_48#_M1005_g N_X_c_619_n 6.66379e-19 $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_193_48#_M1013_g N_X_c_619_n 0.00849619f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_193_48#_M1020_g N_X_c_619_n 3.55395e-19 $X=2.34 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A_193_48#_M1002_g N_X_c_620_n 2.99553e-19 $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A_193_48#_c_160_n X 0.0015671f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_193_48#_c_161_n X 0.0012794f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_193_48#_c_159_n X 0.0177465f $X=2.34 $Y=1.527 $X2=0 $Y2=0
cc_233 N_A_193_48#_c_160_n N_X_c_626_n 0.00942645f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_193_48#_M1002_g N_X_c_622_n 0.00252852f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_193_48#_M1005_g N_X_c_622_n 0.0038796f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_193_48#_c_152_n N_X_c_622_n 0.0253315f $X=2.81 $Y=1.455 $X2=0 $Y2=0
cc_237 N_A_193_48#_c_159_n N_X_c_622_n 0.0134482f $X=2.34 $Y=1.527 $X2=0 $Y2=0
cc_238 N_A_193_48#_c_164_n N_A_892_392#_M1004_d 0.00202164f $X=4.975 $Y=2.125
+ $X2=-0.19 $Y2=-0.245
cc_239 N_A_193_48#_c_164_n N_A_892_392#_c_673_n 0.0179042f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_240 N_A_193_48#_c_207_p N_A_892_392#_c_673_n 0.0172613f $X=5.06 $Y=2.57 $X2=0
+ $Y2=0
cc_241 N_A_193_48#_M1008_d N_A_892_392#_c_669_n 0.00225108f $X=4.91 $Y=1.96
+ $X2=0 $Y2=0
cc_242 N_A_193_48#_c_164_n N_A_892_392#_c_669_n 0.00358435f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_243 N_A_193_48#_c_207_p N_A_892_392#_c_669_n 0.012787f $X=5.06 $Y=2.57 $X2=0
+ $Y2=0
cc_244 N_A_193_48#_c_165_n N_A_892_392#_c_671_n 0.0255098f $X=5.06 $Y=2.3 $X2=0
+ $Y2=0
cc_245 N_A_193_48#_c_207_p N_A_892_392#_c_671_n 0.0283023f $X=5.06 $Y=2.57 $X2=0
+ $Y2=0
cc_246 N_A_193_48#_M1002_g N_VGND_c_700_n 0.0105578f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_193_48#_M1005_g N_VGND_c_700_n 4.79292e-19 $X=1.48 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_193_48#_M1002_g N_VGND_c_701_n 4.62568e-19 $X=1.04 $Y=0.74 $X2=0
+ $Y2=0
cc_249 N_A_193_48#_M1005_g N_VGND_c_701_n 0.00870114f $X=1.48 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A_193_48#_M1013_g N_VGND_c_701_n 0.00167001f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_251 N_A_193_48#_M1013_g N_VGND_c_702_n 6.04497e-19 $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_252 N_A_193_48#_M1020_g N_VGND_c_702_n 0.014379f $X=2.34 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_193_48#_c_152_n N_VGND_c_702_n 0.0214009f $X=2.81 $Y=1.455 $X2=0
+ $Y2=0
cc_254 N_A_193_48#_c_153_n N_VGND_c_702_n 0.0528834f $X=2.895 $Y=1.29 $X2=0
+ $Y2=0
cc_255 N_A_193_48#_c_155_n N_VGND_c_702_n 0.0146661f $X=2.98 $Y=0.34 $X2=0 $Y2=0
cc_256 N_A_193_48#_c_159_n N_VGND_c_702_n 0.00214634f $X=2.34 $Y=1.527 $X2=0
+ $Y2=0
cc_257 N_A_193_48#_c_154_n N_VGND_c_703_n 0.00519468f $X=3.5 $Y=0.34 $X2=0 $Y2=0
cc_258 N_A_193_48#_c_177_p N_VGND_c_703_n 0.00482934f $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_259 N_A_193_48#_M1013_g N_VGND_c_705_n 0.00434272f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_260 N_A_193_48#_M1020_g N_VGND_c_705_n 0.00383152f $X=2.34 $Y=0.74 $X2=0
+ $Y2=0
cc_261 N_A_193_48#_M1002_g N_VGND_c_707_n 0.00429299f $X=1.04 $Y=0.74 $X2=0
+ $Y2=0
cc_262 N_A_193_48#_M1005_g N_VGND_c_707_n 0.00383152f $X=1.48 $Y=0.74 $X2=0
+ $Y2=0
cc_263 N_A_193_48#_c_154_n N_VGND_c_708_n 0.0566428f $X=3.5 $Y=0.34 $X2=0 $Y2=0
cc_264 N_A_193_48#_c_155_n N_VGND_c_708_n 0.0121867f $X=2.98 $Y=0.34 $X2=0 $Y2=0
cc_265 N_A_193_48#_M1002_g N_VGND_c_711_n 0.00847623f $X=1.04 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A_193_48#_M1005_g N_VGND_c_711_n 0.0075764f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_193_48#_M1013_g N_VGND_c_711_n 0.00820284f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_193_48#_M1020_g N_VGND_c_711_n 0.0075754f $X=2.34 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_193_48#_c_154_n N_VGND_c_711_n 0.0322874f $X=3.5 $Y=0.34 $X2=0 $Y2=0
cc_270 N_A_193_48#_c_155_n N_VGND_c_711_n 0.00660921f $X=2.98 $Y=0.34 $X2=0
+ $Y2=0
cc_271 N_A_193_48#_c_153_n N_A_618_94#_c_800_n 0.0262213f $X=2.895 $Y=1.29 $X2=0
+ $Y2=0
cc_272 N_A_193_48#_c_154_n N_A_618_94#_c_800_n 0.0127218f $X=3.5 $Y=0.34 $X2=0
+ $Y2=0
cc_273 N_A_193_48#_M1007_d N_A_618_94#_c_791_n 0.00176461f $X=3.525 $Y=0.47
+ $X2=0 $Y2=0
cc_274 N_A_193_48#_c_154_n N_A_618_94#_c_791_n 0.0042894f $X=3.5 $Y=0.34 $X2=0
+ $Y2=0
cc_275 N_A_193_48#_c_156_n N_A_618_94#_c_791_n 0.03855f $X=3.66 $Y=1.375 $X2=0
+ $Y2=0
cc_276 N_A_193_48#_c_177_p N_A_618_94#_c_791_n 0.0167224f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_277 N_A_193_48#_c_153_n N_A_618_94#_c_792_n 0.0140746f $X=2.895 $Y=1.29 $X2=0
+ $Y2=0
cc_278 N_A_193_48#_c_156_n N_A_618_94#_c_792_n 0.0140592f $X=3.66 $Y=1.375 $X2=0
+ $Y2=0
cc_279 N_A_193_48#_c_164_n N_A_618_94#_c_794_n 0.00468152f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_280 N_A_193_48#_c_164_n N_A_618_94#_c_798_n 0.00590868f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_281 N_A_27_368#_M1019_g N_A1_M1006_g 0.0285527f $X=3.88 $Y=0.79 $X2=0 $Y2=0
cc_282 N_A_27_368#_c_319_n N_A1_c_470_n 0.0223437f $X=3.8 $Y=2.045 $X2=0 $Y2=0
cc_283 N_A_27_368#_M1019_g N_A1_c_470_n 0.0195598f $X=3.88 $Y=0.79 $X2=0 $Y2=0
cc_284 N_A_27_368#_c_317_n N_A1_c_470_n 0.0084556f $X=3.8 $Y=1.837 $X2=0 $Y2=0
cc_285 N_A_27_368#_M1019_g A1 0.00126428f $X=3.88 $Y=0.79 $X2=0 $Y2=0
cc_286 N_A_27_368#_c_331_n N_VPWR_M1016_d 0.0142647f $X=3.15 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_287 N_A_27_368#_c_331_n N_VPWR_M1012_s 0.00392025f $X=3.15 $Y=2.475 $X2=0
+ $Y2=0
cc_288 N_A_27_368#_c_331_n N_VPWR_M1017_s 0.0346593f $X=3.15 $Y=2.475 $X2=0
+ $Y2=0
cc_289 N_A_27_368#_c_322_n N_VPWR_M1017_s 0.00476538f $X=3.235 $Y=2.39 $X2=0
+ $Y2=0
cc_290 N_A_27_368#_c_321_n N_VPWR_c_540_n 0.0103139f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_291 N_A_27_368#_c_331_n N_VPWR_c_540_n 0.0236138f $X=3.15 $Y=2.475 $X2=0
+ $Y2=0
cc_292 N_A_27_368#_c_331_n N_VPWR_c_541_n 0.0166996f $X=3.15 $Y=2.475 $X2=0
+ $Y2=0
cc_293 N_A_27_368#_c_319_n N_VPWR_c_542_n 0.00803176f $X=3.8 $Y=2.045 $X2=0
+ $Y2=0
cc_294 N_A_27_368#_c_321_n N_VPWR_c_545_n 0.0159324f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_295 N_A_27_368#_c_318_n N_VPWR_c_547_n 0.00461464f $X=3.35 $Y=2.045 $X2=0
+ $Y2=0
cc_296 N_A_27_368#_c_319_n N_VPWR_c_547_n 0.00445602f $X=3.8 $Y=2.045 $X2=0
+ $Y2=0
cc_297 N_A_27_368#_c_318_n N_VPWR_c_552_n 0.0111714f $X=3.35 $Y=2.045 $X2=0
+ $Y2=0
cc_298 N_A_27_368#_c_331_n N_VPWR_c_552_n 0.0539598f $X=3.15 $Y=2.475 $X2=0
+ $Y2=0
cc_299 N_A_27_368#_c_318_n N_VPWR_c_539_n 0.00775099f $X=3.35 $Y=2.045 $X2=0
+ $Y2=0
cc_300 N_A_27_368#_c_319_n N_VPWR_c_539_n 0.00858864f $X=3.8 $Y=2.045 $X2=0
+ $Y2=0
cc_301 N_A_27_368#_c_321_n N_VPWR_c_539_n 0.0131546f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_302 N_A_27_368#_c_331_n N_VPWR_c_539_n 0.052919f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_303 N_A_27_368#_c_331_n N_X_M1011_d 0.00549176f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_304 N_A_27_368#_c_331_n N_X_M1014_d 0.00549507f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_305 N_A_27_368#_c_331_n N_X_c_623_n 0.0561701f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_306 N_A_27_368#_c_331_n N_X_c_626_n 0.0137955f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_307 N_A_27_368#_c_323_n N_X_c_626_n 0.0106111f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A_27_368#_c_313_n N_VGND_c_700_n 0.026158f $X=0.31 $Y=0.515 $X2=0 $Y2=0
cc_309 N_A_27_368#_M1007_g N_VGND_c_708_n 7.82275e-19 $X=3.45 $Y=0.79 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_M1019_g N_VGND_c_708_n 0.00435309f $X=3.88 $Y=0.79 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_M1019_g N_VGND_c_711_n 0.00428698f $X=3.88 $Y=0.79 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_c_313_n N_VGND_c_711_n 0.0142062f $X=0.31 $Y=0.515 $X2=0
+ $Y2=0
cc_313 N_A_27_368#_c_313_n N_VGND_c_712_n 0.0172202f $X=0.31 $Y=0.515 $X2=0
+ $Y2=0
cc_314 N_A_27_368#_M1007_g N_A_618_94#_c_791_n 0.0111584f $X=3.45 $Y=0.79 $X2=0
+ $Y2=0
cc_315 N_A_27_368#_M1019_g N_A_618_94#_c_791_n 0.0167517f $X=3.88 $Y=0.79 $X2=0
+ $Y2=0
cc_316 N_A_27_368#_c_317_n N_A_618_94#_c_791_n 2.51936e-19 $X=3.8 $Y=1.837 $X2=0
+ $Y2=0
cc_317 N_A_27_368#_M1019_g N_A_618_94#_c_798_n 0.00501111f $X=3.88 $Y=0.79 $X2=0
+ $Y2=0
cc_318 N_A2_M1003_g N_A1_M1006_g 0.0248487f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_319 N_A2_c_414_n N_A1_c_470_n 0.0343186f $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_320 A2 N_A1_c_470_n 2.60921e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_321 N_A2_c_413_n N_A1_c_470_n 0.0236977f $X=5.285 $Y=1.667 $X2=0 $Y2=0
cc_322 N_A2_M1003_g N_A1_c_471_n 0.00895007f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_323 N_A2_M1009_g N_A1_c_471_n 0.00894529f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_324 N_A2_M1009_g N_A1_c_473_n 0.00674476f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_325 A2 N_A1_c_474_n 0.0255537f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_326 N_A2_c_413_n N_A1_c_474_n 0.0209507f $X=5.285 $Y=1.667 $X2=0 $Y2=0
cc_327 N_A2_c_415_n N_A1_c_479_n 0.00887292f $X=5.285 $Y=1.885 $X2=0 $Y2=0
cc_328 N_A2_M1009_g N_A1_M1010_g 0.0218553f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_329 A2 A1 0.0285452f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_330 N_A2_c_413_n A1 0.00274698f $X=5.285 $Y=1.667 $X2=0 $Y2=0
cc_331 A2 N_VPWR_c_544_n 0.0211423f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_332 N_A2_c_414_n N_VPWR_c_548_n 0.00278257f $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_333 N_A2_c_415_n N_VPWR_c_548_n 0.00278257f $X=5.285 $Y=1.885 $X2=0 $Y2=0
cc_334 N_A2_c_414_n N_VPWR_c_539_n 0.00353905f $X=4.835 $Y=1.885 $X2=0 $Y2=0
cc_335 N_A2_c_415_n N_VPWR_c_539_n 0.00353905f $X=5.285 $Y=1.885 $X2=0 $Y2=0
cc_336 N_A2_c_414_n N_A_892_392#_c_673_n 0.0067586f $X=4.835 $Y=1.885 $X2=0
+ $Y2=0
cc_337 N_A2_c_415_n N_A_892_392#_c_673_n 5.16405e-19 $X=5.285 $Y=1.885 $X2=0
+ $Y2=0
cc_338 N_A2_c_414_n N_A_892_392#_c_669_n 0.00858774f $X=4.835 $Y=1.885 $X2=0
+ $Y2=0
cc_339 N_A2_c_415_n N_A_892_392#_c_669_n 0.0125587f $X=5.285 $Y=1.885 $X2=0
+ $Y2=0
cc_340 N_A2_c_414_n N_A_892_392#_c_670_n 0.0024094f $X=4.835 $Y=1.885 $X2=0
+ $Y2=0
cc_341 N_A2_c_414_n N_A_892_392#_c_671_n 6.77696e-19 $X=4.835 $Y=1.885 $X2=0
+ $Y2=0
cc_342 N_A2_c_415_n N_A_892_392#_c_671_n 0.011216f $X=5.285 $Y=1.885 $X2=0 $Y2=0
cc_343 A2 N_A_892_392#_c_671_n 0.0286493f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_344 N_A2_c_413_n N_A_892_392#_c_671_n 5.15027e-19 $X=5.285 $Y=1.667 $X2=0
+ $Y2=0
cc_345 N_A2_M1003_g N_VGND_c_703_n 0.0017139f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_346 N_A2_M1003_g N_VGND_c_704_n 4.44858e-19 $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_347 N_A2_M1009_g N_VGND_c_704_n 0.00728275f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_348 N_A2_M1003_g N_VGND_c_711_n 9.49986e-19 $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_349 N_A2_M1009_g N_VGND_c_711_n 7.97988e-19 $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_350 N_A2_M1003_g N_A_618_94#_c_793_n 5.46534e-19 $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_351 N_A2_M1003_g N_A_618_94#_c_794_n 0.0118284f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_352 A2 N_A_618_94#_c_794_n 0.00603618f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_353 N_A2_c_413_n N_A_618_94#_c_794_n 0.00183773f $X=5.285 $Y=1.667 $X2=0
+ $Y2=0
cc_354 N_A2_M1003_g N_A_618_94#_c_795_n 0.00720634f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_355 N_A2_M1009_g N_A_618_94#_c_796_n 0.0121607f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_356 A2 N_A_618_94#_c_796_n 0.0742946f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_357 N_A2_M1009_g N_A_618_94#_c_797_n 5.70901e-19 $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_358 N_A2_M1003_g N_A_618_94#_c_799_n 9.00612e-19 $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_359 A2 N_A_618_94#_c_799_n 0.0209604f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_360 N_A2_c_413_n N_A_618_94#_c_799_n 0.00232511f $X=5.285 $Y=1.667 $X2=0
+ $Y2=0
cc_361 N_A1_c_470_n N_VPWR_c_542_n 0.00466147f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_362 N_A1_c_479_n N_VPWR_c_544_n 0.00681294f $X=5.735 $Y=1.885 $X2=0 $Y2=0
cc_363 N_A1_c_470_n N_VPWR_c_548_n 0.0044313f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_364 N_A1_c_479_n N_VPWR_c_548_n 0.0044313f $X=5.735 $Y=1.885 $X2=0 $Y2=0
cc_365 N_A1_c_470_n N_VPWR_c_539_n 0.00853935f $X=4.385 $Y=1.885 $X2=0 $Y2=0
cc_366 N_A1_c_479_n N_VPWR_c_539_n 0.00856939f $X=5.735 $Y=1.885 $X2=0 $Y2=0
cc_367 N_A1_c_470_n N_A_892_392#_c_673_n 0.0052946f $X=4.385 $Y=1.885 $X2=0
+ $Y2=0
cc_368 N_A1_c_479_n N_A_892_392#_c_669_n 0.00332677f $X=5.735 $Y=1.885 $X2=0
+ $Y2=0
cc_369 N_A1_c_470_n N_A_892_392#_c_670_n 0.00383257f $X=4.385 $Y=1.885 $X2=0
+ $Y2=0
cc_370 N_A1_c_479_n N_A_892_392#_c_671_n 0.0110021f $X=5.735 $Y=1.885 $X2=0
+ $Y2=0
cc_371 N_A1_M1006_g N_VGND_c_703_n 0.0104443f $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_372 N_A1_c_471_n N_VGND_c_703_n 0.0190951f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_373 N_A1_c_471_n N_VGND_c_704_n 0.0190272f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_374 N_A1_M1010_g N_VGND_c_704_n 0.012705f $X=5.74 $Y=0.945 $X2=0 $Y2=0
cc_375 N_A1_c_472_n N_VGND_c_708_n 0.00730708f $X=4.455 $Y=0.18 $X2=0 $Y2=0
cc_376 N_A1_c_471_n N_VGND_c_709_n 0.0187698f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_377 N_A1_c_471_n N_VGND_c_710_n 0.00769733f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_378 N_A1_c_471_n N_VGND_c_711_n 0.0364405f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_379 N_A1_c_472_n N_VGND_c_711_n 0.0106516f $X=4.455 $Y=0.18 $X2=0 $Y2=0
cc_380 N_A1_M1006_g N_A_618_94#_c_793_n 0.00490618f $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_381 N_A1_M1006_g N_A_618_94#_c_794_n 0.0120608f $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_382 N_A1_c_470_n N_A_618_94#_c_794_n 0.00116046f $X=4.385 $Y=1.885 $X2=0
+ $Y2=0
cc_383 A1 N_A_618_94#_c_794_n 0.0261629f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_384 N_A1_M1006_g N_A_618_94#_c_795_n 6.06182e-19 $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_385 N_A1_c_471_n N_A_618_94#_c_795_n 0.00449787f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_386 N_A1_c_473_n N_A_618_94#_c_796_n 8.68351e-19 $X=5.735 $Y=1.43 $X2=0 $Y2=0
cc_387 N_A1_M1010_g N_A_618_94#_c_796_n 0.0121208f $X=5.74 $Y=0.945 $X2=0 $Y2=0
cc_388 N_A1_M1010_g N_A_618_94#_c_797_n 0.00753506f $X=5.74 $Y=0.945 $X2=0 $Y2=0
cc_389 N_A1_M1006_g N_A_618_94#_c_798_n 0.00691928f $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_390 N_A1_c_470_n N_A_618_94#_c_798_n 0.00303582f $X=4.385 $Y=1.885 $X2=0
+ $Y2=0
cc_391 A1 N_A_618_94#_c_798_n 0.0128713f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_392 N_VPWR_M1012_s N_X_c_623_n 0.0020349f $X=1.58 $Y=1.84 $X2=0 $Y2=0
cc_393 N_VPWR_c_544_n N_A_892_392#_c_669_n 0.012272f $X=5.96 $Y=2.115 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_548_n N_A_892_392#_c_669_n 0.0594312f $X=5.875 $Y=3.33 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_539_n N_A_892_392#_c_669_n 0.0328875f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_396 N_VPWR_c_542_n N_A_892_392#_c_670_n 0.0119239f $X=4.11 $Y=2.635 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_548_n N_A_892_392#_c_670_n 0.0233459f $X=5.875 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_539_n N_A_892_392#_c_670_n 0.0126535f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_399 N_VPWR_c_544_n N_A_892_392#_c_671_n 0.0640156f $X=5.96 $Y=2.115 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_544_n N_A_618_94#_c_796_n 3.21367e-19 $X=5.96 $Y=2.115 $X2=0
+ $Y2=0
cc_401 N_X_c_618_n N_VGND_M1005_d 0.00176461f $X=1.96 $Y=1.035 $X2=0 $Y2=0
cc_402 N_X_c_617_n N_VGND_c_700_n 0.0232433f $X=1.255 $Y=0.515 $X2=0 $Y2=0
cc_403 N_X_c_617_n N_VGND_c_701_n 0.0288482f $X=1.255 $Y=0.515 $X2=0 $Y2=0
cc_404 N_X_c_618_n N_VGND_c_701_n 0.0153337f $X=1.96 $Y=1.035 $X2=0 $Y2=0
cc_405 N_X_c_619_n N_VGND_c_701_n 0.0154978f $X=2.125 $Y=0.515 $X2=0 $Y2=0
cc_406 N_X_c_618_n N_VGND_c_702_n 0.00626822f $X=1.96 $Y=1.035 $X2=0 $Y2=0
cc_407 N_X_c_619_n N_VGND_c_702_n 0.021337f $X=2.125 $Y=0.515 $X2=0 $Y2=0
cc_408 N_X_c_619_n N_VGND_c_705_n 0.0109942f $X=2.125 $Y=0.515 $X2=0 $Y2=0
cc_409 N_X_c_617_n N_VGND_c_707_n 0.00861184f $X=1.255 $Y=0.515 $X2=0 $Y2=0
cc_410 N_X_c_617_n N_VGND_c_711_n 0.00712813f $X=1.255 $Y=0.515 $X2=0 $Y2=0
cc_411 N_X_c_619_n N_VGND_c_711_n 0.00904371f $X=2.125 $Y=0.515 $X2=0 $Y2=0
cc_412 N_VGND_c_703_n N_A_618_94#_c_793_n 0.013328f $X=4.665 $Y=0.77 $X2=0 $Y2=0
cc_413 N_VGND_c_708_n N_A_618_94#_c_793_n 0.00670736f $X=4.5 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_711_n N_A_618_94#_c_793_n 0.0100487f $X=6 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_M1006_s N_A_618_94#_c_794_n 0.00250873f $X=4.455 $Y=0.625 $X2=0
+ $Y2=0
cc_416 N_VGND_c_703_n N_A_618_94#_c_794_n 0.0192006f $X=4.665 $Y=0.77 $X2=0
+ $Y2=0
cc_417 N_VGND_c_703_n N_A_618_94#_c_795_n 0.0122347f $X=4.665 $Y=0.77 $X2=0
+ $Y2=0
cc_418 N_VGND_c_704_n N_A_618_94#_c_795_n 0.0122347f $X=5.525 $Y=0.77 $X2=0
+ $Y2=0
cc_419 N_VGND_c_709_n N_A_618_94#_c_795_n 0.00528395f $X=5.36 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_711_n N_A_618_94#_c_795_n 0.00668313f $X=6 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_M1009_d N_A_618_94#_c_796_n 0.00176461f $X=5.385 $Y=0.625 $X2=0
+ $Y2=0
cc_422 N_VGND_c_704_n N_A_618_94#_c_796_n 0.0152916f $X=5.525 $Y=0.77 $X2=0
+ $Y2=0
cc_423 N_VGND_c_704_n N_A_618_94#_c_797_n 0.0127625f $X=5.525 $Y=0.77 $X2=0
+ $Y2=0
cc_424 N_VGND_c_710_n N_A_618_94#_c_797_n 0.00712528f $X=6 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_711_n N_A_618_94#_c_797_n 0.0102037f $X=6 $Y=0 $X2=0 $Y2=0
