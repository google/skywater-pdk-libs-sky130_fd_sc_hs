* File: sky130_fd_sc_hs__a31oi_4.spice
* Created: Tue Sep  1 19:53:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a31oi_4.pex.spice"
.subckt sky130_fd_sc_hs__a31oi_4  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 N_A_30_74#_M1005_d N_A3_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1007 N_A_30_74#_M1007_d N_A3_M1007_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1028 N_A_30_74#_M1007_d N_A3_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1029 N_A_30_74#_M1029_d N_A3_M1029_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_475_74#_M1001_d N_A2_M1001_g N_A_30_74#_M1029_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1004 N_A_475_74#_M1001_d N_A2_M1004_g N_A_30_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_475_74#_M1008_d N_A2_M1008_g N_A_30_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1023 N_A_475_74#_M1008_d N_A2_M1023_g N_A_30_74#_M1023_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.202325 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75003.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g N_A_475_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.19805 AS=0.2109 PD=2.07 PS=1.31 NRD=0.804 NRS=23.508 M=1 R=4.93333
+ SA=75000.2 SB=75003.6 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A1_M1002_g N_A_475_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=1.31 NRD=0 NRS=23.508 M=1 R=4.93333 SA=75000.9
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1002_d N_A1_M1012_g N_A_475_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1017 N_Y_M1017_d N_A1_M1017_g N_A_475_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1017_d N_B1_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.40885 PD=1.09 PS=1.845 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1027 N_Y_M1027_d N_B1_M1027_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.40885 PD=2.05 PS=1.845 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_368#_M1006_d N_A3_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007.8 A=0.168 P=2.54 MULT=1
MM1010 N_A_27_368#_M1010_d N_A3_M1010_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75007.4 A=0.168 P=2.54 MULT=1
MM1011 N_A_27_368#_M1010_d N_A3_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75006.9 A=0.168 P=2.54 MULT=1
MM1013 N_A_27_368#_M1013_d N_A3_M1013_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75006.5 A=0.168 P=2.54 MULT=1
MM1014 N_A_27_368#_M1013_d N_A2_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75006 A=0.168 P=2.54 MULT=1
MM1018 N_A_27_368#_M1018_d N_A2_M1018_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.5 SB=75005.5 A=0.168 P=2.54 MULT=1
MM1020 N_A_27_368#_M1018_d N_A2_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003 SB=75005.1 A=0.168 P=2.54 MULT=1
MM1021 N_A_27_368#_M1021_d N_A2_M1021_g N_VPWR_M1020_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75004.6 A=0.168 P=2.54 MULT=1
MM1015 N_A_27_368#_M1021_d N_A1_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004 SB=75004.1 A=0.168 P=2.54 MULT=1
MM1016 N_A_27_368#_M1016_d N_A1_M1016_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1.12
+ AD=0.4648 AS=0.196 PD=1.95 PS=1.47 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1019 N_A_27_368#_M1016_d N_A1_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1.12
+ AD=0.4648 AS=0.224 PD=1.95 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75005.4 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1024 N_A_27_368#_M1024_d N_A1_M1024_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1848 AS=0.224 PD=1.45 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75006 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_27_368#_M1024_d VPB PSHORT L=0.15 W=1.12
+ AD=0.1792 AS=0.1848 PD=1.44 PS=1.45 NRD=5.2599 NRS=7.0329 M=1 R=7.46667
+ SA=75006.5 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1022 N_Y_M1003_d N_B1_M1022_g N_A_27_368#_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1792 AS=0.168 PD=1.44 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.9 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1025 N_Y_M1025_d N_B1_M1025_g N_A_27_368#_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1026 N_Y_M1025_d N_B1_M1026_g N_A_27_368#_M1026_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX30_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_hs__a31oi_4.pxi.spice"
*
.ends
*
*
