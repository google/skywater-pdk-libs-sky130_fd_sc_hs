* File: sky130_fd_sc_hs__mux2_4.pxi.spice
* Created: Tue Sep  1 20:07:47 2020
* 
x_PM_SKY130_FD_SC_HS__MUX2_4%S N_S_c_158_n N_S_M1016_g N_S_M1003_g N_S_M1001_g
+ N_S_c_167_n N_S_M1002_g N_S_M1024_g N_S_c_168_n N_S_M1007_g N_S_c_169_n
+ N_S_c_178_p N_S_c_179_p N_S_c_184_p N_S_c_170_n N_S_c_162_n N_S_c_163_n
+ N_S_c_185_p S N_S_c_164_n N_S_c_165_n PM_SKY130_FD_SC_HS__MUX2_4%S
x_PM_SKY130_FD_SC_HS__MUX2_4%A_27_368# N_A_27_368#_M1003_s N_A_27_368#_M1016_s
+ N_A_27_368#_c_303_n N_A_27_368#_M1000_g N_A_27_368#_M1005_g
+ N_A_27_368#_M1010_g N_A_27_368#_c_304_n N_A_27_368#_M1020_g
+ N_A_27_368#_c_305_n N_A_27_368#_c_317_n N_A_27_368#_c_306_n
+ N_A_27_368#_c_322_n N_A_27_368#_c_326_n N_A_27_368#_c_307_n
+ N_A_27_368#_c_308_n N_A_27_368#_c_309_n N_A_27_368#_c_298_n
+ N_A_27_368#_c_299_n N_A_27_368#_c_300_n N_A_27_368#_c_311_n
+ N_A_27_368#_c_301_n N_A_27_368#_c_354_n N_A_27_368#_c_302_n
+ PM_SKY130_FD_SC_HS__MUX2_4%A_27_368#
x_PM_SKY130_FD_SC_HS__MUX2_4%A_193_241# N_A_193_241#_M1017_s
+ N_A_193_241#_M1022_s N_A_193_241#_M1025_d N_A_193_241#_M1004_s
+ N_A_193_241#_M1008_s N_A_193_241#_M1019_s N_A_193_241#_c_433_n
+ N_A_193_241#_c_466_n N_A_193_241#_M1006_g N_A_193_241#_M1009_g
+ N_A_193_241#_c_435_n N_A_193_241#_c_436_n N_A_193_241#_c_437_n
+ N_A_193_241#_c_438_n N_A_193_241#_c_468_n N_A_193_241#_M1011_g
+ N_A_193_241#_M1014_g N_A_193_241#_c_440_n N_A_193_241#_M1021_g
+ N_A_193_241#_c_442_n N_A_193_241#_c_443_n N_A_193_241#_c_470_n
+ N_A_193_241#_M1012_g N_A_193_241#_c_444_n N_A_193_241#_M1023_g
+ N_A_193_241#_c_446_n N_A_193_241#_c_447_n N_A_193_241#_c_448_n
+ N_A_193_241#_c_472_n N_A_193_241#_M1013_g N_A_193_241#_c_449_n
+ N_A_193_241#_c_450_n N_A_193_241#_c_451_n N_A_193_241#_c_452_n
+ N_A_193_241#_c_453_n N_A_193_241#_c_454_n N_A_193_241#_c_455_n
+ N_A_193_241#_c_475_n N_A_193_241#_c_476_n N_A_193_241#_c_477_n
+ N_A_193_241#_c_456_n N_A_193_241#_c_537_p N_A_193_241#_c_457_n
+ N_A_193_241#_c_458_n N_A_193_241#_c_478_n N_A_193_241#_c_459_n
+ N_A_193_241#_c_460_n N_A_193_241#_c_461_n N_A_193_241#_c_462_n
+ N_A_193_241#_c_463_n N_A_193_241#_c_480_n N_A_193_241#_c_464_n
+ PM_SKY130_FD_SC_HS__MUX2_4%A_193_241#
x_PM_SKY130_FD_SC_HS__MUX2_4%A0 N_A0_M1017_g N_A0_c_667_n N_A0_M1004_g
+ N_A0_M1022_g N_A0_c_668_n N_A0_M1008_g A0 N_A0_c_666_n
+ PM_SKY130_FD_SC_HS__MUX2_4%A0
x_PM_SKY130_FD_SC_HS__MUX2_4%A1 N_A1_c_713_n N_A1_M1018_g N_A1_M1015_g
+ N_A1_c_714_n N_A1_M1019_g N_A1_M1025_g A1 A1 N_A1_c_711_n N_A1_c_712_n
+ PM_SKY130_FD_SC_HS__MUX2_4%A1
x_PM_SKY130_FD_SC_HS__MUX2_4%VPWR N_VPWR_M1016_d N_VPWR_M1011_d N_VPWR_M1013_d
+ N_VPWR_M1007_s N_VPWR_M1020_d N_VPWR_c_757_n N_VPWR_c_758_n N_VPWR_c_759_n
+ N_VPWR_c_760_n N_VPWR_c_761_n N_VPWR_c_762_n N_VPWR_c_763_n N_VPWR_c_764_n
+ N_VPWR_c_765_n N_VPWR_c_766_n N_VPWR_c_767_n VPWR N_VPWR_c_768_n
+ N_VPWR_c_769_n N_VPWR_c_756_n N_VPWR_c_771_n N_VPWR_c_772_n
+ PM_SKY130_FD_SC_HS__MUX2_4%VPWR
x_PM_SKY130_FD_SC_HS__MUX2_4%X N_X_M1009_d N_X_M1021_d N_X_M1006_s N_X_M1012_s
+ N_X_c_857_n N_X_c_858_n N_X_c_859_n N_X_c_860_n X X X N_X_c_861_n X
+ PM_SKY130_FD_SC_HS__MUX2_4%X
x_PM_SKY130_FD_SC_HS__MUX2_4%A_722_391# N_A_722_391#_M1002_d
+ N_A_722_391#_M1004_d N_A_722_391#_c_921_n N_A_722_391#_c_922_n
+ N_A_722_391#_c_923_n N_A_722_391#_c_924_n
+ PM_SKY130_FD_SC_HS__MUX2_4%A_722_391#
x_PM_SKY130_FD_SC_HS__MUX2_4%A_936_391# N_A_936_391#_M1000_s
+ N_A_936_391#_M1018_d N_A_936_391#_c_970_n N_A_936_391#_c_971_n
+ N_A_936_391#_c_972_n N_A_936_391#_c_973_n N_A_936_391#_c_974_n
+ PM_SKY130_FD_SC_HS__MUX2_4%A_936_391#
x_PM_SKY130_FD_SC_HS__MUX2_4%VGND N_VGND_M1003_d N_VGND_M1014_s N_VGND_M1023_s
+ N_VGND_M1024_s N_VGND_M1010_s N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n
+ N_VGND_c_1019_n N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n
+ N_VGND_c_1023_n N_VGND_c_1024_n N_VGND_c_1025_n VGND N_VGND_c_1026_n
+ N_VGND_c_1027_n N_VGND_c_1028_n N_VGND_c_1029_n N_VGND_c_1030_n
+ N_VGND_c_1031_n N_VGND_c_1032_n PM_SKY130_FD_SC_HS__MUX2_4%VGND
x_PM_SKY130_FD_SC_HS__MUX2_4%A_709_119# N_A_709_119#_M1001_d
+ N_A_709_119#_M1015_s N_A_709_119#_c_1122_n N_A_709_119#_c_1123_n
+ N_A_709_119#_c_1124_n N_A_709_119#_c_1125_n N_A_709_119#_c_1126_n
+ N_A_709_119#_c_1127_n PM_SKY130_FD_SC_HS__MUX2_4%A_709_119#
x_PM_SKY130_FD_SC_HS__MUX2_4%A_937_119# N_A_937_119#_M1005_d
+ N_A_937_119#_M1017_d N_A_937_119#_c_1182_n N_A_937_119#_c_1183_n
+ N_A_937_119#_c_1188_n N_A_937_119#_c_1184_n N_A_937_119#_c_1199_n
+ PM_SKY130_FD_SC_HS__MUX2_4%A_937_119#
cc_1 VNB N_S_c_158_n 0.0270854f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_S_M1003_g 0.0294058f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.81
cc_3 VNB N_S_M1001_g 0.0228248f $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=0.915
cc_4 VNB N_S_M1024_g 0.0216899f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.915
cc_5 VNB N_S_c_162_n 0.00152914f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=1.6
cc_6 VNB N_S_c_163_n 0.00633555f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.6
cc_7 VNB N_S_c_164_n 0.00610825f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_8 VNB N_S_c_165_n 0.0276622f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=1.657
cc_9 VNB N_A_27_368#_M1005_g 0.0215488f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=1.88
cc_10 VNB N_A_27_368#_M1010_g 0.0232446f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.915
cc_11 VNB N_A_27_368#_c_298_n 3.75525e-19 $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.135
cc_12 VNB N_A_27_368#_c_299_n 0.00212795f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.24
cc_13 VNB N_A_27_368#_c_300_n 0.0447788f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_14 VNB N_A_27_368#_c_301_n 0.0242993f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.657
cc_15 VNB N_A_27_368#_c_302_n 0.0355754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_193_241#_c_433_n 0.00622475f $X=-0.19 $Y=-0.245 $X2=3.985
+ $Y2=2.455
cc_17 VNB N_A_193_241#_M1009_g 0.0119056f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.24
cc_18 VNB N_A_193_241#_c_435_n 0.0188836f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.765
cc_19 VNB N_A_193_241#_c_436_n 0.0125025f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=2.155
cc_20 VNB N_A_193_241#_c_437_n 0.00590914f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=1.6
cc_21 VNB N_A_193_241#_c_438_n 0.0126506f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.6
cc_22 VNB N_A_193_241#_M1014_g 0.011601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_193_241#_c_440_n 0.0274798f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_24 VNB N_A_193_241#_M1021_g 0.0112763f $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=1.657
cc_25 VNB N_A_193_241#_c_442_n 0.00575392f $X=-0.19 $Y=-0.245 $X2=3.535
+ $Y2=1.657
cc_26 VNB N_A_193_241#_c_443_n 0.0149832f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.657
cc_27 VNB N_A_193_241#_c_444_n 0.016028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_193_241#_M1023_g 0.0129289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_193_241#_c_446_n 0.219476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_193_241#_c_447_n 0.0261311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_193_241#_c_448_n 0.00887312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_193_241#_c_449_n 0.0853864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_193_241#_c_450_n 0.0201574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_193_241#_c_451_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_193_241#_c_452_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_193_241#_c_453_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_193_241#_c_454_n 0.00467671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_193_241#_c_455_n 0.0313614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_193_241#_c_456_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_193_241#_c_457_n 0.012433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_193_241#_c_458_n 0.0165854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_193_241#_c_459_n 0.0302575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_193_241#_c_460_n 0.00938153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_193_241#_c_461_n 0.00139572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_193_241#_c_462_n 0.0022133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_193_241#_c_463_n 0.0133735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_193_241#_c_464_n 0.0171429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A0_M1017_g 0.0448307f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_49 VNB N_A0_M1022_g 0.0336114f $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=0.915
cc_50 VNB N_A0_c_666_n 0.0250441f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.78
cc_51 VNB N_A1_M1015_g 0.0337961f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.81
cc_52 VNB N_A1_M1025_g 0.0391319f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=2.455
cc_53 VNB N_A1_c_711_n 0.00508237f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.05
cc_54 VNB N_A1_c_712_n 0.0281232f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.135
cc_55 VNB N_VPWR_c_756_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_X_c_857_n 0.00243486f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=2.455
cc_57 VNB N_X_c_858_n 0.00541625f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=1.435
cc_58 VNB N_X_c_859_n 7.61737e-19 $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.915
cc_59 VNB N_X_c_860_n 0.00215099f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.88
cc_60 VNB N_X_c_861_n 0.00882506f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=1.6
cc_61 VNB N_VGND_c_1016_n 0.0228137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1017_n 0.00298812f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.78
cc_63 VNB N_VGND_c_1018_n 0.0157969f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=2.24
cc_64 VNB N_VGND_c_1019_n 0.0205418f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=1.6
cc_65 VNB N_VGND_c_1020_n 0.0195912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1021_n 0.0128294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1022_n 0.0234806f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_68 VNB N_VGND_c_1023_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_69 VNB N_VGND_c_1024_n 0.0190194f $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=1.657
cc_70 VNB N_VGND_c_1025_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=1.657
cc_71 VNB N_VGND_c_1026_n 0.0196457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1027_n 0.0171982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1028_n 0.0724602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1029_n 0.434755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1030_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1031_n 0.00625894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1032_n 0.00536684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_709_119#_c_1122_n 0.00267057f $X=-0.19 $Y=-0.245 $X2=3.47
+ $Y2=0.915
cc_79 VNB N_A_709_119#_c_1123_n 0.00289807f $X=-0.19 $Y=-0.245 $X2=3.535
+ $Y2=1.88
cc_80 VNB N_A_709_119#_c_1124_n 0.0407711f $X=-0.19 $Y=-0.245 $X2=3.535
+ $Y2=2.455
cc_81 VNB N_A_709_119#_c_1125_n 0.00218005f $X=-0.19 $Y=-0.245 $X2=3.97
+ $Y2=0.915
cc_82 VNB N_A_709_119#_c_1126_n 0.00740417f $X=-0.19 $Y=-0.245 $X2=3.985
+ $Y2=1.88
cc_83 VNB N_A_709_119#_c_1127_n 0.00609138f $X=-0.19 $Y=-0.245 $X2=3.985
+ $Y2=2.455
cc_84 VNB N_A_937_119#_c_1182_n 0.00160098f $X=-0.19 $Y=-0.245 $X2=3.47
+ $Y2=0.915
cc_85 VNB N_A_937_119#_c_1183_n 0.00224578f $X=-0.19 $Y=-0.245 $X2=3.535
+ $Y2=1.88
cc_86 VNB N_A_937_119#_c_1184_n 0.00151525f $X=-0.19 $Y=-0.245 $X2=3.97
+ $Y2=0.915
cc_87 VPB N_S_c_158_n 0.031122f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_88 VPB N_S_c_167_n 0.016863f $X=-0.19 $Y=1.66 $X2=3.535 $Y2=1.88
cc_89 VPB N_S_c_168_n 0.016456f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=1.88
cc_90 VPB N_S_c_169_n 8.63879e-19 $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.05
cc_91 VPB N_S_c_170_n 0.00123359f $X=-0.19 $Y=1.66 $X2=3.08 $Y2=2.155
cc_92 VPB N_S_c_163_n 0.00697023f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_93 VPB N_S_c_164_n 0.00234496f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_94 VPB N_S_c_165_n 0.0334557f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=1.657
cc_95 VPB N_A_27_368#_c_303_n 0.0170611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_368#_c_304_n 0.0178255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_368#_c_305_n 0.0101859f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.135
cc_98 VPB N_A_27_368#_c_306_n 0.022783f $X=-0.19 $Y=1.66 $X2=2.995 $Y2=2.24
cc_99 VPB N_A_27_368#_c_307_n 0.00263937f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_100 VPB N_A_27_368#_c_308_n 0.00109397f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_101 VPB N_A_27_368#_c_309_n 0.0020303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_368#_c_299_n 0.00390775f $X=-0.19 $Y=1.66 $X2=1.59 $Y2=2.24
cc_103 VPB N_A_27_368#_c_311_n 0.00710642f $X=-0.19 $Y=1.66 $X2=3.535 $Y2=1.657
cc_104 VPB N_A_27_368#_c_301_n 0.0127137f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.657
cc_105 VPB N_A_27_368#_c_302_n 0.0438388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_193_241#_c_433_n 0.0110376f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=2.455
cc_107 VPB N_A_193_241#_c_466_n 0.0242848f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=2.455
cc_108 VPB N_A_193_241#_c_438_n 0.00873592f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_109 VPB N_A_193_241#_c_468_n 0.0233074f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_110 VPB N_A_193_241#_c_443_n 0.00559939f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.657
cc_111 VPB N_A_193_241#_c_470_n 0.023312f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=1.657
cc_112 VPB N_A_193_241#_c_448_n 0.00369733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_193_241#_c_472_n 0.0244274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_193_241#_c_454_n 0.00179237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_193_241#_c_455_n 0.0266663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_193_241#_c_475_n 0.00738474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_193_241#_c_476_n 0.0105261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_193_241#_c_477_n 0.00724744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_193_241#_c_478_n 0.0327264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_193_241#_c_459_n 0.0139269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_193_241#_c_480_n 0.0169392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_193_241#_c_464_n 0.017241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A0_c_667_n 0.0192231f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.81
cc_124 VPB N_A0_c_668_n 0.0159235f $X=-0.19 $Y=1.66 $X2=3.535 $Y2=1.88
cc_125 VPB N_A0_c_666_n 0.0326337f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.78
cc_126 VPB N_A1_c_713_n 0.0159386f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_127 VPB N_A1_c_714_n 0.0203775f $X=-0.19 $Y=1.66 $X2=3.47 $Y2=1.435
cc_128 VPB N_A1_c_711_n 0.00361007f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.05
cc_129 VPB N_A1_c_712_n 0.0345759f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.135
cc_130 VPB N_VPWR_c_757_n 0.0112079f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=2.455
cc_131 VPB N_VPWR_c_758_n 0.00802818f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.135
cc_132 VPB N_VPWR_c_759_n 0.00802264f $X=-0.19 $Y=1.66 $X2=3.08 $Y2=1.765
cc_133 VPB N_VPWR_c_760_n 0.00870426f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_134 VPB N_VPWR_c_761_n 0.00687743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_762_n 0.0232884f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_136 VPB N_VPWR_c_763_n 0.00631622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_764_n 0.0203178f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_138 VPB N_VPWR_c_765_n 0.00631953f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_139 VPB N_VPWR_c_766_n 0.0207444f $X=-0.19 $Y=1.66 $X2=3.535 $Y2=1.657
cc_140 VPB N_VPWR_c_767_n 0.00478125f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.657
cc_141 VPB N_VPWR_c_768_n 0.025094f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.78
cc_142 VPB N_VPWR_c_769_n 0.0862348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_756_n 0.0986956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_771_n 0.0270295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_772_n 0.00631622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_X_c_857_n 5.32607e-19 $X=-0.19 $Y=1.66 $X2=3.535 $Y2=2.455
cc_147 VPB N_X_c_859_n 0.00278809f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=0.915
cc_148 VPB N_X_c_861_n 7.84116e-19 $X=-0.19 $Y=1.66 $X2=3.165 $Y2=1.6
cc_149 VPB N_A_722_391#_c_921_n 0.00357339f $X=-0.19 $Y=1.66 $X2=3.47 $Y2=0.915
cc_150 VPB N_A_722_391#_c_922_n 0.0214742f $X=-0.19 $Y=1.66 $X2=3.535 $Y2=2.455
cc_151 VPB N_A_722_391#_c_923_n 0.00220397f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=0.915
cc_152 VPB N_A_722_391#_c_924_n 0.0177469f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=0.915
cc_153 VPB N_A_936_391#_c_970_n 0.0116889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_936_391#_c_971_n 0.00548534f $X=-0.19 $Y=1.66 $X2=3.47 $Y2=0.915
cc_155 VPB N_A_936_391#_c_972_n 0.00261476f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=0.915
cc_156 VPB N_A_936_391#_c_973_n 0.0162879f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=0.915
cc_157 VPB N_A_936_391#_c_974_n 0.00256835f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.78
cc_158 N_S_c_168_n N_A_27_368#_c_303_n 0.0267268f $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_159 N_S_M1024_g N_A_27_368#_M1005_g 0.0210679f $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_160 N_S_c_158_n N_A_27_368#_c_305_n 0.00589403f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_161 N_S_c_158_n N_A_27_368#_c_317_n 0.0111908f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_162 N_S_c_178_p N_A_27_368#_c_317_n 0.0165225f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_163 N_S_c_179_p N_A_27_368#_c_317_n 0.0137412f $X=0.835 $Y=2.135 $X2=0 $Y2=0
cc_164 N_S_c_164_n N_A_27_368#_c_317_n 0.00532192f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_165 N_S_c_158_n N_A_27_368#_c_306_n 0.00780197f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_166 N_S_c_167_n N_A_27_368#_c_322_n 0.00585856f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_167 N_S_c_178_p N_A_27_368#_c_322_n 0.00866703f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_168 N_S_c_184_p N_A_27_368#_c_322_n 0.086688f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_169 N_S_c_185_p N_A_27_368#_c_322_n 0.00803741f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_170 N_S_c_167_n N_A_27_368#_c_326_n 0.00978564f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_171 N_S_c_168_n N_A_27_368#_c_326_n 7.88787e-19 $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_172 N_S_c_184_p N_A_27_368#_c_326_n 0.0138308f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_173 N_S_c_170_n N_A_27_368#_c_326_n 0.003559f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_174 N_S_c_167_n N_A_27_368#_c_307_n 0.00974419f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_175 N_S_c_168_n N_A_27_368#_c_307_n 0.00865897f $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_176 N_S_c_163_n N_A_27_368#_c_307_n 0.0176104f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_177 N_S_c_165_n N_A_27_368#_c_307_n 0.0081812f $X=3.97 $Y=1.657 $X2=0 $Y2=0
cc_178 N_S_c_167_n N_A_27_368#_c_308_n 0.00315153f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_179 N_S_c_170_n N_A_27_368#_c_308_n 0.0138662f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_180 N_S_c_163_n N_A_27_368#_c_308_n 0.0143813f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_181 N_S_c_165_n N_A_27_368#_c_308_n 0.00183128f $X=3.97 $Y=1.657 $X2=0 $Y2=0
cc_182 N_S_c_167_n N_A_27_368#_c_309_n 3.29415e-19 $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_183 N_S_c_168_n N_A_27_368#_c_309_n 0.0018024f $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_184 N_S_c_165_n N_A_27_368#_c_309_n 0.00490257f $X=3.97 $Y=1.657 $X2=0 $Y2=0
cc_185 N_S_c_163_n N_A_27_368#_c_298_n 0.0277655f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_186 N_S_c_165_n N_A_27_368#_c_298_n 0.0150349f $X=3.97 $Y=1.657 $X2=0 $Y2=0
cc_187 N_S_c_158_n N_A_27_368#_c_300_n 0.00161792f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_188 N_S_M1003_g N_A_27_368#_c_300_n 0.00855288f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_189 N_S_c_164_n N_A_27_368#_c_300_n 0.013094f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_190 N_S_c_158_n N_A_27_368#_c_311_n 0.00211987f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_191 N_S_c_169_n N_A_27_368#_c_311_n 0.00606518f $X=0.75 $Y=2.05 $X2=0 $Y2=0
cc_192 N_S_c_179_p N_A_27_368#_c_311_n 0.0115465f $X=0.835 $Y=2.135 $X2=0 $Y2=0
cc_193 N_S_c_164_n N_A_27_368#_c_311_n 0.00127779f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_194 N_S_c_158_n N_A_27_368#_c_301_n 0.0119239f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_195 N_S_M1003_g N_A_27_368#_c_301_n 0.00436189f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_196 N_S_c_169_n N_A_27_368#_c_301_n 0.00470158f $X=0.75 $Y=2.05 $X2=0 $Y2=0
cc_197 N_S_c_164_n N_A_27_368#_c_301_n 0.0329253f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_198 N_S_c_178_p N_A_27_368#_c_354_n 0.0111307f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_199 N_S_c_165_n N_A_27_368#_c_302_n 0.0209787f $X=3.97 $Y=1.657 $X2=0 $Y2=0
cc_200 N_S_c_158_n N_A_193_241#_c_466_n 0.0285902f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_201 N_S_c_178_p N_A_193_241#_c_466_n 0.0144382f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_202 N_S_c_185_p N_A_193_241#_c_466_n 0.00199304f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_203 N_S_c_164_n N_A_193_241#_c_466_n 0.00475287f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_204 N_S_M1003_g N_A_193_241#_M1009_g 0.0166337f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_205 N_S_c_178_p N_A_193_241#_c_468_n 3.83075e-19 $X=1.505 $Y=2.135 $X2=0
+ $Y2=0
cc_206 N_S_c_184_p N_A_193_241#_c_468_n 0.00698328f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_207 N_S_c_185_p N_A_193_241#_c_468_n 0.00888333f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_208 N_S_c_162_n N_A_193_241#_c_443_n 2.07238e-19 $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_209 N_S_c_184_p N_A_193_241#_c_470_n 0.0129318f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_210 N_S_c_185_p N_A_193_241#_c_470_n 6.00352e-19 $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_211 N_S_M1001_g N_A_193_241#_M1023_g 0.00801147f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_212 N_S_M1001_g N_A_193_241#_c_446_n 0.0103003f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_213 N_S_M1024_g N_A_193_241#_c_446_n 0.0103107f $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_214 N_S_M1001_g N_A_193_241#_c_447_n 0.00702575f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_215 N_S_c_184_p N_A_193_241#_c_447_n 0.00104864f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_216 N_S_c_162_n N_A_193_241#_c_447_n 9.10335e-19 $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_217 N_S_c_162_n N_A_193_241#_c_448_n 0.00573519f $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_218 N_S_c_165_n N_A_193_241#_c_448_n 0.00702575f $X=3.97 $Y=1.657 $X2=0 $Y2=0
cc_219 N_S_c_167_n N_A_193_241#_c_472_n 0.0243198f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_220 N_S_c_184_p N_A_193_241#_c_472_n 0.0159472f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_221 N_S_c_170_n N_A_193_241#_c_472_n 0.00307514f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_222 N_S_c_162_n N_A_193_241#_c_472_n 0.00261042f $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_223 N_S_c_165_n N_A_193_241#_c_472_n 0.0020534f $X=3.97 $Y=1.657 $X2=0 $Y2=0
cc_224 N_S_c_158_n N_A_193_241#_c_450_n 0.0196188f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_225 N_S_M1003_g N_A_193_241#_c_450_n 0.00854554f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_226 N_S_c_164_n N_A_193_241#_c_450_n 0.00313316f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_227 N_S_c_169_n N_VPWR_M1016_d 0.00530254f $X=0.75 $Y=2.05 $X2=-0.19
+ $Y2=-0.245
cc_228 N_S_c_178_p N_VPWR_M1016_d 0.00424661f $X=1.505 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_229 N_S_c_179_p N_VPWR_M1016_d 0.00468788f $X=0.835 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_230 N_S_c_184_p N_VPWR_M1011_d 0.00953446f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_231 N_S_c_184_p N_VPWR_M1013_d 0.00285122f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_232 N_S_c_170_n N_VPWR_M1013_d 0.00332957f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_233 N_S_c_158_n N_VPWR_c_757_n 0.00432031f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_234 N_S_c_167_n N_VPWR_c_759_n 0.00475883f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_235 N_S_c_168_n N_VPWR_c_760_n 0.00518461f $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_236 N_S_c_167_n N_VPWR_c_764_n 0.00418024f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_237 N_S_c_168_n N_VPWR_c_764_n 0.00329149f $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_238 N_S_c_158_n N_VPWR_c_756_n 0.00508379f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_239 N_S_c_167_n N_VPWR_c_756_n 0.00544287f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_240 N_S_c_168_n N_VPWR_c_756_n 0.00544287f $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_241 N_S_c_158_n N_VPWR_c_771_n 0.00481134f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_242 N_S_c_178_p N_X_M1006_s 0.00854178f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_243 N_S_c_185_p N_X_M1006_s 0.00260597f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_244 N_S_c_184_p N_X_M1012_s 0.00863676f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_245 N_S_c_158_n N_X_c_857_n 3.60404e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_246 N_S_c_178_p N_X_c_857_n 0.0289881f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_247 N_S_c_185_p N_X_c_857_n 0.00629455f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_248 N_S_c_164_n N_X_c_857_n 0.032f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_249 N_S_c_164_n N_X_c_858_n 8.05573e-19 $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_250 N_S_M1001_g N_X_c_859_n 2.44849e-19 $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_251 N_S_c_184_p N_X_c_859_n 0.0295758f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_252 N_S_c_170_n N_X_c_859_n 0.0100274f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_253 N_S_c_162_n N_X_c_859_n 0.0226861f $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_254 N_S_M1001_g N_X_c_860_n 0.00101895f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_255 N_S_c_184_p N_X_c_861_n 0.029062f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_256 N_S_c_185_p N_X_c_861_n 0.00257766f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_257 N_S_c_168_n N_A_722_391#_c_921_n 0.0108466f $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_258 N_S_c_167_n N_A_722_391#_c_923_n 0.00453579f $X=3.535 $Y=1.88 $X2=0 $Y2=0
cc_259 N_S_c_168_n N_A_722_391#_c_923_n 0.00929261f $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_260 N_S_c_168_n N_A_936_391#_c_972_n 8.53536e-19 $X=3.985 $Y=1.88 $X2=0 $Y2=0
cc_261 N_S_M1003_g N_VGND_c_1016_n 0.0074703f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_262 N_S_c_164_n N_VGND_c_1016_n 0.00525943f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_263 N_S_M1001_g N_VGND_c_1018_n 0.0108034f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_264 N_S_c_162_n N_VGND_c_1018_n 0.0152459f $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_265 N_S_c_163_n N_VGND_c_1018_n 0.00752017f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_266 N_S_M1001_g N_VGND_c_1020_n 6.03908e-19 $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_267 N_S_M1024_g N_VGND_c_1020_n 0.0133679f $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_268 N_S_M1003_g N_VGND_c_1022_n 0.00473385f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_269 N_S_M1003_g N_VGND_c_1029_n 0.00508379f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_270 N_S_M1001_g N_VGND_c_1029_n 9.39239e-19 $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_271 N_S_M1024_g N_VGND_c_1029_n 7.88961e-19 $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_272 N_S_M1001_g N_A_709_119#_c_1122_n 0.00735844f $X=3.47 $Y=0.915 $X2=0
+ $Y2=0
cc_273 N_S_M1024_g N_A_709_119#_c_1122_n 0.00277359f $X=3.97 $Y=0.915 $X2=0
+ $Y2=0
cc_274 N_S_M1001_g N_A_709_119#_c_1123_n 0.00334323f $X=3.47 $Y=0.915 $X2=0
+ $Y2=0
cc_275 N_S_c_163_n N_A_709_119#_c_1123_n 0.0188868f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_276 N_S_c_165_n N_A_709_119#_c_1123_n 0.0043641f $X=3.97 $Y=1.657 $X2=0 $Y2=0
cc_277 N_S_M1024_g N_A_709_119#_c_1126_n 0.0157322f $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_278 N_S_c_165_n N_A_709_119#_c_1126_n 2.09528e-19 $X=3.97 $Y=1.657 $X2=0
+ $Y2=0
cc_279 N_S_M1024_g N_A_937_119#_c_1183_n 2.92953e-19 $X=3.97 $Y=0.915 $X2=0
+ $Y2=0
cc_280 N_A_27_368#_c_305_n N_A_193_241#_c_466_n 7.7052e-19 $X=0.265 $Y=2.39
+ $X2=0 $Y2=0
cc_281 N_A_27_368#_c_317_n N_A_193_241#_c_466_n 0.0114142f $X=1.165 $Y=2.475
+ $X2=0 $Y2=0
cc_282 N_A_27_368#_c_306_n N_A_193_241#_c_466_n 5.08122e-19 $X=0.445 $Y=2.475
+ $X2=0 $Y2=0
cc_283 N_A_27_368#_c_322_n N_A_193_241#_c_468_n 0.0129745f $X=3.335 $Y=2.58
+ $X2=0 $Y2=0
cc_284 N_A_27_368#_c_354_n N_A_193_241#_c_468_n 0.0023078f $X=1.25 $Y=2.475
+ $X2=0 $Y2=0
cc_285 N_A_27_368#_c_322_n N_A_193_241#_c_470_n 0.0136487f $X=3.335 $Y=2.58
+ $X2=0 $Y2=0
cc_286 N_A_27_368#_M1005_g N_A_193_241#_c_446_n 0.0103003f $X=4.61 $Y=0.915
+ $X2=0 $Y2=0
cc_287 N_A_27_368#_M1010_g N_A_193_241#_c_446_n 0.00991298f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_288 N_A_27_368#_c_322_n N_A_193_241#_c_472_n 0.0135726f $X=3.335 $Y=2.58
+ $X2=0 $Y2=0
cc_289 N_A_27_368#_c_326_n N_A_193_241#_c_472_n 0.00357033f $X=3.42 $Y=2.495
+ $X2=0 $Y2=0
cc_290 N_A_27_368#_M1010_g N_A_193_241#_c_449_n 0.0193743f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_291 N_A_27_368#_c_299_n N_A_193_241#_c_454_n 0.0132241f $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_292 N_A_27_368#_c_302_n N_A_193_241#_c_454_n 0.00154688f $X=5.04 $Y=1.657
+ $X2=0 $Y2=0
cc_293 N_A_27_368#_c_299_n N_A_193_241#_c_464_n 3.11698e-19 $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_294 N_A_27_368#_c_302_n N_A_193_241#_c_464_n 0.0187061f $X=5.04 $Y=1.657
+ $X2=0 $Y2=0
cc_295 N_A_27_368#_c_317_n N_VPWR_M1016_d 0.00675622f $X=1.165 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_296 N_A_27_368#_c_322_n N_VPWR_M1011_d 0.00865418f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_297 N_A_27_368#_c_322_n N_VPWR_M1013_d 0.0125765f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_298 N_A_27_368#_c_326_n N_VPWR_M1013_d 0.00420304f $X=3.42 $Y=2.495 $X2=0
+ $Y2=0
cc_299 N_A_27_368#_c_308_n N_VPWR_M1013_d 0.00139828f $X=3.505 $Y=2.02 $X2=0
+ $Y2=0
cc_300 N_A_27_368#_c_317_n N_VPWR_c_757_n 0.0225065f $X=1.165 $Y=2.475 $X2=0
+ $Y2=0
cc_301 N_A_27_368#_c_306_n N_VPWR_c_757_n 0.0088922f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_302 N_A_27_368#_c_322_n N_VPWR_c_758_n 0.0252358f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_303 N_A_27_368#_c_322_n N_VPWR_c_759_n 0.0256372f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_304 N_A_27_368#_c_303_n N_VPWR_c_760_n 0.00894559f $X=4.605 $Y=1.88 $X2=0
+ $Y2=0
cc_305 N_A_27_368#_c_304_n N_VPWR_c_761_n 0.0123918f $X=5.055 $Y=1.88 $X2=0
+ $Y2=0
cc_306 N_A_27_368#_c_322_n N_VPWR_c_762_n 0.00692546f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_307 N_A_27_368#_c_354_n N_VPWR_c_762_n 0.00268263f $X=1.25 $Y=2.475 $X2=0
+ $Y2=0
cc_308 N_A_27_368#_c_322_n N_VPWR_c_764_n 0.00149698f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_c_303_n N_VPWR_c_766_n 0.00332316f $X=4.605 $Y=1.88 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_c_304_n N_VPWR_c_766_n 0.00332316f $X=5.055 $Y=1.88 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_c_322_n N_VPWR_c_768_n 0.0128691f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_c_303_n N_VPWR_c_756_n 0.00544287f $X=4.605 $Y=1.88 $X2=0
+ $Y2=0
cc_313 N_A_27_368#_c_304_n N_VPWR_c_756_n 0.00544287f $X=5.055 $Y=1.88 $X2=0
+ $Y2=0
cc_314 N_A_27_368#_c_317_n N_VPWR_c_756_n 0.0136101f $X=1.165 $Y=2.475 $X2=0
+ $Y2=0
cc_315 N_A_27_368#_c_306_n N_VPWR_c_756_n 0.0122756f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_316 N_A_27_368#_c_322_n N_VPWR_c_756_n 0.0428516f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_317 N_A_27_368#_c_354_n N_VPWR_c_756_n 0.00478779f $X=1.25 $Y=2.475 $X2=0
+ $Y2=0
cc_318 N_A_27_368#_c_306_n N_VPWR_c_771_n 0.0107406f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_319 N_A_27_368#_c_322_n N_X_M1006_s 0.00755126f $X=3.335 $Y=2.58 $X2=0 $Y2=0
cc_320 N_A_27_368#_c_354_n N_X_M1006_s 0.00638397f $X=1.25 $Y=2.475 $X2=0 $Y2=0
cc_321 N_A_27_368#_c_322_n N_X_M1012_s 0.0112288f $X=3.335 $Y=2.58 $X2=0 $Y2=0
cc_322 N_A_27_368#_c_307_n N_A_722_391#_M1002_d 0.00219742f $X=3.915 $Y=2.02
+ $X2=-0.19 $Y2=-0.245
cc_323 N_A_27_368#_c_303_n N_A_722_391#_c_921_n 0.015091f $X=4.605 $Y=1.88 $X2=0
+ $Y2=0
cc_324 N_A_27_368#_c_304_n N_A_722_391#_c_921_n 0.0139612f $X=5.055 $Y=1.88
+ $X2=0 $Y2=0
cc_325 N_A_27_368#_c_307_n N_A_722_391#_c_921_n 0.0060041f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_326 N_A_27_368#_c_299_n N_A_722_391#_c_921_n 0.0138858f $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_327 N_A_27_368#_c_302_n N_A_722_391#_c_921_n 0.00290564f $X=5.04 $Y=1.657
+ $X2=0 $Y2=0
cc_328 N_A_27_368#_c_303_n N_A_722_391#_c_923_n 0.00148763f $X=4.605 $Y=1.88
+ $X2=0 $Y2=0
cc_329 N_A_27_368#_c_322_n N_A_722_391#_c_923_n 0.0144217f $X=3.335 $Y=2.58
+ $X2=0 $Y2=0
cc_330 N_A_27_368#_c_326_n N_A_722_391#_c_923_n 0.0163401f $X=3.42 $Y=2.495
+ $X2=0 $Y2=0
cc_331 N_A_27_368#_c_307_n N_A_722_391#_c_923_n 0.0156265f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_332 N_A_27_368#_c_304_n N_A_722_391#_c_924_n 0.00483173f $X=5.055 $Y=1.88
+ $X2=0 $Y2=0
cc_333 N_A_27_368#_c_303_n N_A_936_391#_c_972_n 0.00728288f $X=4.605 $Y=1.88
+ $X2=0 $Y2=0
cc_334 N_A_27_368#_c_304_n N_A_936_391#_c_972_n 0.0175583f $X=5.055 $Y=1.88
+ $X2=0 $Y2=0
cc_335 N_A_27_368#_c_307_n N_A_936_391#_c_972_n 0.00281087f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_336 N_A_27_368#_c_299_n N_A_936_391#_c_972_n 0.0252424f $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_337 N_A_27_368#_c_302_n N_A_936_391#_c_972_n 0.0080882f $X=5.04 $Y=1.657
+ $X2=0 $Y2=0
cc_338 N_A_27_368#_c_300_n N_VGND_c_1016_n 0.0288933f $X=0.435 $Y=0.635 $X2=0
+ $Y2=0
cc_339 N_A_27_368#_M1005_g N_VGND_c_1020_n 0.00585775f $X=4.61 $Y=0.915 $X2=0
+ $Y2=0
cc_340 N_A_27_368#_M1010_g N_VGND_c_1021_n 0.00351782f $X=5.04 $Y=0.915 $X2=0
+ $Y2=0
cc_341 N_A_27_368#_c_300_n N_VGND_c_1022_n 0.0153192f $X=0.435 $Y=0.635 $X2=0
+ $Y2=0
cc_342 N_A_27_368#_M1005_g N_VGND_c_1029_n 9.39239e-19 $X=4.61 $Y=0.915 $X2=0
+ $Y2=0
cc_343 N_A_27_368#_M1010_g N_VGND_c_1029_n 9.39239e-19 $X=5.04 $Y=0.915 $X2=0
+ $Y2=0
cc_344 N_A_27_368#_c_300_n N_VGND_c_1029_n 0.0175003f $X=0.435 $Y=0.635 $X2=0
+ $Y2=0
cc_345 N_A_27_368#_c_307_n N_A_709_119#_c_1123_n 0.00335306f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_346 N_A_27_368#_M1005_g N_A_709_119#_c_1126_n 0.0150485f $X=4.61 $Y=0.915
+ $X2=0 $Y2=0
cc_347 N_A_27_368#_M1010_g N_A_709_119#_c_1126_n 0.0133803f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_348 N_A_27_368#_c_307_n N_A_709_119#_c_1126_n 0.00174523f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_349 N_A_27_368#_c_298_n N_A_709_119#_c_1126_n 0.0131287f $X=4.085 $Y=1.6
+ $X2=0 $Y2=0
cc_350 N_A_27_368#_c_299_n N_A_709_119#_c_1126_n 0.0679154f $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_302_n N_A_709_119#_c_1126_n 0.00816766f $X=5.04 $Y=1.657
+ $X2=0 $Y2=0
cc_352 N_A_27_368#_M1010_g N_A_709_119#_c_1127_n 4.91777e-19 $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_353 N_A_27_368#_M1005_g N_A_937_119#_c_1183_n 0.00472551f $X=4.61 $Y=0.915
+ $X2=0 $Y2=0
cc_354 N_A_27_368#_M1010_g N_A_937_119#_c_1183_n 0.00553184f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_355 N_A_27_368#_M1010_g N_A_937_119#_c_1188_n 0.0101743f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_356 N_A_27_368#_M1010_g N_A_937_119#_c_1184_n 3.25189e-19 $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_357 N_A_193_241#_c_456_n N_A0_M1017_g 0.0121398f $X=7.26 $Y=0.34 $X2=0 $Y2=0
cc_358 N_A_193_241#_c_475_n N_A0_c_667_n 0.00216762f $X=6.385 $Y=1.95 $X2=0
+ $Y2=0
cc_359 N_A_193_241#_c_476_n N_A0_c_667_n 0.0109486f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_360 N_A_193_241#_c_456_n N_A0_M1022_g 0.013161f $X=7.26 $Y=0.34 $X2=0 $Y2=0
cc_361 N_A_193_241#_c_476_n N_A0_c_668_n 0.0131287f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_362 N_A_193_241#_c_454_n A0 0.02833f $X=6.3 $Y=1.615 $X2=0 $Y2=0
cc_363 N_A_193_241#_c_455_n A0 3.51297e-19 $X=6.23 $Y=1.615 $X2=0 $Y2=0
cc_364 N_A_193_241#_c_476_n A0 0.0330885f $X=8.195 $Y=2.075 $X2=0 $Y2=0
cc_365 N_A_193_241#_c_454_n N_A0_c_666_n 0.00239229f $X=6.3 $Y=1.615 $X2=0 $Y2=0
cc_366 N_A_193_241#_c_455_n N_A0_c_666_n 0.0182643f $X=6.23 $Y=1.615 $X2=0 $Y2=0
cc_367 N_A_193_241#_c_475_n N_A0_c_666_n 0.00367265f $X=6.385 $Y=1.95 $X2=0
+ $Y2=0
cc_368 N_A_193_241#_c_476_n N_A0_c_666_n 0.00870706f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_369 N_A_193_241#_c_476_n N_A1_c_713_n 0.0108827f $X=8.195 $Y=2.075 $X2=-0.19
+ $Y2=-0.245
cc_370 N_A_193_241#_c_537_p N_A1_M1015_g 0.00708055f $X=7.425 $Y=0.495 $X2=0
+ $Y2=0
cc_371 N_A_193_241#_c_457_n N_A1_M1015_g 0.0102487f $X=8.19 $Y=0.34 $X2=0 $Y2=0
cc_372 N_A_193_241#_c_462_n N_A1_M1015_g 0.00203192f $X=7.425 $Y=0.34 $X2=0
+ $Y2=0
cc_373 N_A_193_241#_c_476_n N_A1_c_714_n 0.0204034f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_374 N_A_193_241#_c_478_n N_A1_c_714_n 0.0153381f $X=8.36 $Y=2.465 $X2=0 $Y2=0
cc_375 N_A_193_241#_c_459_n N_A1_c_714_n 4.83444e-19 $X=8.44 $Y=1.95 $X2=0 $Y2=0
cc_376 N_A_193_241#_c_537_p N_A1_M1025_g 6.1326e-19 $X=7.425 $Y=0.495 $X2=0
+ $Y2=0
cc_377 N_A_193_241#_c_457_n N_A1_M1025_g 0.0142468f $X=8.19 $Y=0.34 $X2=0 $Y2=0
cc_378 N_A_193_241#_c_459_n N_A1_M1025_g 0.00991507f $X=8.44 $Y=1.95 $X2=0 $Y2=0
cc_379 N_A_193_241#_c_463_n N_A1_M1025_g 4.67633e-19 $X=8.357 $Y=1.03 $X2=0
+ $Y2=0
cc_380 N_A_193_241#_c_476_n N_A1_c_711_n 0.0653717f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_381 N_A_193_241#_c_459_n N_A1_c_711_n 0.025097f $X=8.44 $Y=1.95 $X2=0 $Y2=0
cc_382 N_A_193_241#_c_476_n N_A1_c_712_n 0.00932519f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_383 N_A_193_241#_c_459_n N_A1_c_712_n 0.00592795f $X=8.44 $Y=1.95 $X2=0 $Y2=0
cc_384 N_A_193_241#_c_466_n N_VPWR_c_757_n 0.01045f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_385 N_A_193_241#_c_468_n N_VPWR_c_757_n 0.00158022f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_386 N_A_193_241#_c_468_n N_VPWR_c_758_n 0.0073295f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_387 N_A_193_241#_c_470_n N_VPWR_c_758_n 0.0073295f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_388 N_A_193_241#_c_472_n N_VPWR_c_759_n 0.00738277f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_A_193_241#_c_466_n N_VPWR_c_762_n 0.00413917f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_390 N_A_193_241#_c_468_n N_VPWR_c_762_n 0.003294f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_391 N_A_193_241#_c_470_n N_VPWR_c_768_n 0.003294f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_392 N_A_193_241#_c_472_n N_VPWR_c_768_n 0.003294f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_393 N_A_193_241#_c_478_n N_VPWR_c_769_n 0.0146357f $X=8.36 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A_193_241#_c_466_n N_VPWR_c_756_n 0.00400044f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_395 N_A_193_241#_c_468_n N_VPWR_c_756_n 0.00423545f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_396 N_A_193_241#_c_470_n N_VPWR_c_756_n 0.00423545f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_397 N_A_193_241#_c_472_n N_VPWR_c_756_n 0.00426944f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_398 N_A_193_241#_c_478_n N_VPWR_c_756_n 0.0121141f $X=8.36 $Y=2.465 $X2=0
+ $Y2=0
cc_399 N_A_193_241#_c_433_n N_X_c_857_n 0.0118288f $X=1.055 $Y=1.675 $X2=0 $Y2=0
cc_400 N_A_193_241#_c_466_n N_X_c_857_n 0.00732875f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_401 N_A_193_241#_c_438_n N_X_c_857_n 0.00665574f $X=1.675 $Y=1.675 $X2=0
+ $Y2=0
cc_402 N_A_193_241#_c_468_n N_X_c_857_n 0.00521068f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_403 N_A_193_241#_c_450_n N_X_c_857_n 0.00827407f $X=1.22 $Y=1.28 $X2=0 $Y2=0
cc_404 N_A_193_241#_M1009_g N_X_c_858_n 0.00662985f $X=1.22 $Y=0.76 $X2=0 $Y2=0
cc_405 N_A_193_241#_c_435_n N_X_c_858_n 0.00327521f $X=1.615 $Y=0.18 $X2=0 $Y2=0
cc_406 N_A_193_241#_c_437_n N_X_c_858_n 0.00379227f $X=1.675 $Y=1.295 $X2=0
+ $Y2=0
cc_407 N_A_193_241#_c_438_n N_X_c_858_n 0.00250774f $X=1.675 $Y=1.675 $X2=0
+ $Y2=0
cc_408 N_A_193_241#_M1014_g N_X_c_858_n 0.0120726f $X=1.69 $Y=0.76 $X2=0 $Y2=0
cc_409 N_A_193_241#_M1021_g N_X_c_858_n 0.00149354f $X=2.28 $Y=0.76 $X2=0 $Y2=0
cc_410 N_A_193_241#_c_443_n N_X_c_859_n 0.0056737f $X=2.295 $Y=1.675 $X2=0 $Y2=0
cc_411 N_A_193_241#_c_470_n N_X_c_859_n 0.0080241f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_412 N_A_193_241#_c_447_n N_X_c_859_n 0.00715706f $X=2.915 $Y=1.46 $X2=0 $Y2=0
cc_413 N_A_193_241#_c_448_n N_X_c_859_n 0.00282915f $X=2.915 $Y=1.675 $X2=0
+ $Y2=0
cc_414 N_A_193_241#_c_472_n N_X_c_859_n 0.00299757f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_A_193_241#_M1014_g N_X_c_860_n 0.00150338f $X=1.69 $Y=0.76 $X2=0 $Y2=0
cc_416 N_A_193_241#_M1021_g N_X_c_860_n 0.0125712f $X=2.28 $Y=0.76 $X2=0 $Y2=0
cc_417 N_A_193_241#_c_442_n N_X_c_860_n 0.0038955f $X=2.295 $Y=1.295 $X2=0 $Y2=0
cc_418 N_A_193_241#_c_443_n N_X_c_860_n 0.00255008f $X=2.295 $Y=1.675 $X2=0
+ $Y2=0
cc_419 N_A_193_241#_c_444_n N_X_c_860_n 0.00233944f $X=2.635 $Y=0.18 $X2=0 $Y2=0
cc_420 N_A_193_241#_M1023_g N_X_c_860_n 0.021545f $X=2.71 $Y=0.76 $X2=0 $Y2=0
cc_421 N_A_193_241#_c_447_n N_X_c_860_n 0.00253386f $X=2.915 $Y=1.46 $X2=0 $Y2=0
cc_422 N_A_193_241#_c_438_n N_X_c_861_n 0.0148285f $X=1.675 $Y=1.675 $X2=0 $Y2=0
cc_423 N_A_193_241#_c_468_n N_X_c_861_n 0.00779845f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_A_193_241#_c_443_n N_X_c_861_n 0.0148285f $X=2.295 $Y=1.675 $X2=0 $Y2=0
cc_425 N_A_193_241#_c_470_n N_X_c_861_n 0.00795893f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_A_193_241#_c_476_n N_A_722_391#_M1004_d 0.00200574f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_427 N_A_193_241#_M1004_s N_A_722_391#_c_922_n 0.00501822f $X=6.32 $Y=1.96
+ $X2=0 $Y2=0
cc_428 N_A_193_241#_c_476_n N_A_936_391#_M1018_d 0.00200085f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_429 N_A_193_241#_c_454_n N_A_936_391#_c_970_n 0.0270752f $X=6.3 $Y=1.615
+ $X2=0 $Y2=0
cc_430 N_A_193_241#_c_464_n N_A_936_391#_c_970_n 0.0121277f $X=5.78 $Y=1.615
+ $X2=0 $Y2=0
cc_431 N_A_193_241#_M1004_s N_A_936_391#_c_971_n 0.00708736f $X=6.32 $Y=1.96
+ $X2=0 $Y2=0
cc_432 N_A_193_241#_M1008_s N_A_936_391#_c_971_n 0.00585944f $X=7.25 $Y=1.96
+ $X2=0 $Y2=0
cc_433 N_A_193_241#_c_454_n N_A_936_391#_c_971_n 0.00496304f $X=6.3 $Y=1.615
+ $X2=0 $Y2=0
cc_434 N_A_193_241#_c_455_n N_A_936_391#_c_971_n 0.00303812f $X=6.23 $Y=1.615
+ $X2=0 $Y2=0
cc_435 N_A_193_241#_c_476_n N_A_936_391#_c_971_n 0.0679747f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_436 N_A_193_241#_c_477_n N_A_936_391#_c_971_n 0.013893f $X=6.47 $Y=2.075
+ $X2=0 $Y2=0
cc_437 N_A_193_241#_c_454_n N_A_936_391#_c_973_n 0.00864147f $X=6.3 $Y=1.615
+ $X2=0 $Y2=0
cc_438 N_A_193_241#_c_455_n N_A_936_391#_c_973_n 0.00352482f $X=6.23 $Y=1.615
+ $X2=0 $Y2=0
cc_439 N_A_193_241#_c_477_n N_A_936_391#_c_973_n 0.0088683f $X=6.47 $Y=2.075
+ $X2=0 $Y2=0
cc_440 N_A_193_241#_c_476_n N_A_936_391#_c_974_n 0.0176481f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_441 N_A_193_241#_c_478_n N_A_936_391#_c_974_n 0.0172628f $X=8.36 $Y=2.465
+ $X2=0 $Y2=0
cc_442 N_A_193_241#_c_436_n N_VGND_c_1016_n 0.0155675f $X=1.295 $Y=0.18 $X2=0
+ $Y2=0
cc_443 N_A_193_241#_c_450_n N_VGND_c_1016_n 0.0070114f $X=1.22 $Y=1.28 $X2=0
+ $Y2=0
cc_444 N_A_193_241#_M1014_g N_VGND_c_1017_n 0.00786117f $X=1.69 $Y=0.76 $X2=0
+ $Y2=0
cc_445 N_A_193_241#_c_440_n N_VGND_c_1017_n 0.0244461f $X=2.205 $Y=0.18 $X2=0
+ $Y2=0
cc_446 N_A_193_241#_M1021_g N_VGND_c_1017_n 0.00999417f $X=2.28 $Y=0.76 $X2=0
+ $Y2=0
cc_447 N_A_193_241#_M1021_g N_VGND_c_1018_n 0.00138461f $X=2.28 $Y=0.76 $X2=0
+ $Y2=0
cc_448 N_A_193_241#_M1023_g N_VGND_c_1018_n 0.0100627f $X=2.71 $Y=0.76 $X2=0
+ $Y2=0
cc_449 N_A_193_241#_c_446_n N_VGND_c_1018_n 0.0261591f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_450 N_A_193_241#_c_447_n N_VGND_c_1018_n 0.00405865f $X=2.915 $Y=1.46 $X2=0
+ $Y2=0
cc_451 N_A_193_241#_c_446_n N_VGND_c_1019_n 0.0232603f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_452 N_A_193_241#_c_446_n N_VGND_c_1020_n 0.0334796f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_453 N_A_193_241#_c_446_n N_VGND_c_1021_n 0.0277529f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_454 N_A_193_241#_c_449_n N_VGND_c_1021_n 0.00432999f $X=5.705 $Y=1.45 $X2=0
+ $Y2=0
cc_455 N_A_193_241#_c_460_n N_VGND_c_1021_n 0.021907f $X=6.425 $Y=0.515 $X2=0
+ $Y2=0
cc_456 N_A_193_241#_c_436_n N_VGND_c_1024_n 0.0208701f $X=1.295 $Y=0.18 $X2=0
+ $Y2=0
cc_457 N_A_193_241#_c_440_n N_VGND_c_1026_n 0.0241797f $X=2.205 $Y=0.18 $X2=0
+ $Y2=0
cc_458 N_A_193_241#_c_446_n N_VGND_c_1027_n 0.0185474f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_459 N_A_193_241#_c_446_n N_VGND_c_1028_n 0.00710974f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_460 N_A_193_241#_c_457_n N_VGND_c_1028_n 0.0618101f $X=8.19 $Y=0.34 $X2=0
+ $Y2=0
cc_461 N_A_193_241#_c_460_n N_VGND_c_1028_n 0.0933251f $X=6.425 $Y=0.515 $X2=0
+ $Y2=0
cc_462 N_A_193_241#_c_462_n N_VGND_c_1028_n 0.0235818f $X=7.425 $Y=0.34 $X2=0
+ $Y2=0
cc_463 N_A_193_241#_c_435_n N_VGND_c_1029_n 0.00836613f $X=1.615 $Y=0.18 $X2=0
+ $Y2=0
cc_464 N_A_193_241#_c_436_n N_VGND_c_1029_n 0.0114564f $X=1.295 $Y=0.18 $X2=0
+ $Y2=0
cc_465 N_A_193_241#_c_440_n N_VGND_c_1029_n 0.00646961f $X=2.205 $Y=0.18 $X2=0
+ $Y2=0
cc_466 N_A_193_241#_c_444_n N_VGND_c_1029_n 0.00686833f $X=2.635 $Y=0.18 $X2=0
+ $Y2=0
cc_467 N_A_193_241#_c_446_n N_VGND_c_1029_n 0.0624474f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_468 N_A_193_241#_c_451_n N_VGND_c_1029_n 0.00824287f $X=1.69 $Y=0.18 $X2=0
+ $Y2=0
cc_469 N_A_193_241#_c_452_n N_VGND_c_1029_n 0.00829753f $X=2.28 $Y=0.18 $X2=0
+ $Y2=0
cc_470 N_A_193_241#_c_453_n N_VGND_c_1029_n 0.00491962f $X=2.71 $Y=0.18 $X2=0
+ $Y2=0
cc_471 N_A_193_241#_c_457_n N_VGND_c_1029_n 0.0343238f $X=8.19 $Y=0.34 $X2=0
+ $Y2=0
cc_472 N_A_193_241#_c_460_n N_VGND_c_1029_n 0.052653f $X=6.425 $Y=0.515 $X2=0
+ $Y2=0
cc_473 N_A_193_241#_c_462_n N_VGND_c_1029_n 0.0127177f $X=7.425 $Y=0.34 $X2=0
+ $Y2=0
cc_474 N_A_193_241#_c_457_n N_A_709_119#_M1015_s 0.00208352f $X=8.19 $Y=0.34
+ $X2=0 $Y2=0
cc_475 N_A_193_241#_c_446_n N_A_709_119#_c_1122_n 0.00622628f $X=5.63 $Y=0.18
+ $X2=0 $Y2=0
cc_476 N_A_193_241#_c_449_n N_A_709_119#_c_1124_n 0.0135146f $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_477 N_A_193_241#_c_454_n N_A_709_119#_c_1124_n 0.0820582f $X=6.3 $Y=1.615
+ $X2=0 $Y2=0
cc_478 N_A_193_241#_c_455_n N_A_709_119#_c_1124_n 0.0123082f $X=6.23 $Y=1.615
+ $X2=0 $Y2=0
cc_479 N_A_193_241#_c_476_n N_A_709_119#_c_1124_n 0.0113132f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_480 N_A_193_241#_c_537_p N_A_709_119#_c_1124_n 0.0229858f $X=7.425 $Y=0.495
+ $X2=0 $Y2=0
cc_481 N_A_193_241#_c_459_n N_A_709_119#_c_1124_n 0.00893256f $X=8.44 $Y=1.95
+ $X2=0 $Y2=0
cc_482 N_A_193_241#_c_464_n N_A_709_119#_c_1124_n 0.00549303f $X=5.78 $Y=1.615
+ $X2=0 $Y2=0
cc_483 N_A_193_241#_c_457_n N_A_709_119#_c_1125_n 0.0149266f $X=8.19 $Y=0.34
+ $X2=0 $Y2=0
cc_484 N_A_193_241#_c_459_n N_A_709_119#_c_1125_n 0.00142601f $X=8.44 $Y=1.95
+ $X2=0 $Y2=0
cc_485 N_A_193_241#_c_463_n N_A_709_119#_c_1125_n 0.00155021f $X=8.357 $Y=1.03
+ $X2=0 $Y2=0
cc_486 N_A_193_241#_c_449_n N_A_709_119#_c_1127_n 3.54931e-19 $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_487 N_A_193_241#_c_456_n N_A_937_119#_M1017_d 0.00197722f $X=7.26 $Y=0.34
+ $X2=0 $Y2=0
cc_488 N_A_193_241#_M1017_s N_A_937_119#_c_1182_n 0.019235f $X=5.855 $Y=0.37
+ $X2=0 $Y2=0
cc_489 N_A_193_241#_c_449_n N_A_937_119#_c_1182_n 0.009911f $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_490 N_A_193_241#_c_456_n N_A_937_119#_c_1182_n 0.00418581f $X=7.26 $Y=0.34
+ $X2=0 $Y2=0
cc_491 N_A_193_241#_c_460_n N_A_937_119#_c_1182_n 0.0552517f $X=6.425 $Y=0.515
+ $X2=0 $Y2=0
cc_492 N_A_193_241#_c_446_n N_A_937_119#_c_1183_n 0.00557458f $X=5.63 $Y=0.18
+ $X2=0 $Y2=0
cc_493 N_A_193_241#_c_449_n N_A_937_119#_c_1183_n 8.19579e-19 $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_494 N_A_193_241#_c_446_n N_A_937_119#_c_1188_n 0.00156495f $X=5.63 $Y=0.18
+ $X2=0 $Y2=0
cc_495 N_A_193_241#_c_449_n N_A_937_119#_c_1184_n 0.0057997f $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_496 N_A_193_241#_c_456_n N_A_937_119#_c_1199_n 0.0152769f $X=7.26 $Y=0.34
+ $X2=0 $Y2=0
cc_497 N_A0_c_668_n N_A1_c_713_n 0.034704f $X=7.175 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_498 N_A0_M1022_g N_A1_M1015_g 0.022348f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_499 A0 N_A1_c_711_n 0.0211953f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_500 N_A0_c_666_n N_A1_c_711_n 0.0034029f $X=7.16 $Y=1.667 $X2=0 $Y2=0
cc_501 A0 N_A1_c_712_n 2.45568e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_502 N_A0_c_666_n N_A1_c_712_n 0.0223794f $X=7.16 $Y=1.667 $X2=0 $Y2=0
cc_503 N_A0_c_667_n N_VPWR_c_769_n 0.00291649f $X=6.725 $Y=1.885 $X2=0 $Y2=0
cc_504 N_A0_c_668_n N_VPWR_c_769_n 0.00444483f $X=7.175 $Y=1.885 $X2=0 $Y2=0
cc_505 N_A0_c_667_n N_VPWR_c_756_n 0.00364317f $X=6.725 $Y=1.885 $X2=0 $Y2=0
cc_506 N_A0_c_668_n N_VPWR_c_756_n 0.00443368f $X=7.175 $Y=1.885 $X2=0 $Y2=0
cc_507 N_A0_c_667_n N_A_722_391#_c_922_n 0.0140124f $X=6.725 $Y=1.885 $X2=0
+ $Y2=0
cc_508 N_A0_c_668_n N_A_722_391#_c_922_n 0.00533934f $X=7.175 $Y=1.885 $X2=0
+ $Y2=0
cc_509 N_A0_c_667_n N_A_936_391#_c_971_n 0.0124098f $X=6.725 $Y=1.885 $X2=0
+ $Y2=0
cc_510 N_A0_c_668_n N_A_936_391#_c_971_n 0.0118516f $X=7.175 $Y=1.885 $X2=0
+ $Y2=0
cc_511 N_A0_c_667_n N_A_936_391#_c_973_n 0.00314988f $X=6.725 $Y=1.885 $X2=0
+ $Y2=0
cc_512 N_A0_c_668_n N_A_936_391#_c_974_n 0.00160701f $X=7.175 $Y=1.885 $X2=0
+ $Y2=0
cc_513 N_A0_M1017_g N_VGND_c_1028_n 0.00278271f $X=6.71 $Y=0.69 $X2=0 $Y2=0
cc_514 N_A0_M1022_g N_VGND_c_1028_n 0.00278271f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_515 N_A0_M1017_g N_VGND_c_1029_n 0.00357715f $X=6.71 $Y=0.69 $X2=0 $Y2=0
cc_516 N_A0_M1022_g N_VGND_c_1029_n 0.00350534f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_517 N_A0_M1017_g N_A_709_119#_c_1124_n 0.0127036f $X=6.71 $Y=0.69 $X2=0 $Y2=0
cc_518 N_A0_M1022_g N_A_709_119#_c_1124_n 0.0174943f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_519 A0 N_A_709_119#_c_1124_n 0.032153f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_520 N_A0_c_666_n N_A_709_119#_c_1124_n 0.00341313f $X=7.16 $Y=1.667 $X2=0
+ $Y2=0
cc_521 N_A0_M1017_g N_A_937_119#_c_1182_n 0.0112042f $X=6.71 $Y=0.69 $X2=0 $Y2=0
cc_522 N_A0_M1017_g N_A_937_119#_c_1199_n 0.00916617f $X=6.71 $Y=0.69 $X2=0
+ $Y2=0
cc_523 N_A0_M1022_g N_A_937_119#_c_1199_n 0.0030388f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_524 N_A1_c_713_n N_VPWR_c_769_n 0.00445602f $X=7.635 $Y=1.885 $X2=0 $Y2=0
cc_525 N_A1_c_714_n N_VPWR_c_769_n 0.00445602f $X=8.085 $Y=1.885 $X2=0 $Y2=0
cc_526 N_A1_c_713_n N_VPWR_c_756_n 0.00442412f $X=7.635 $Y=1.885 $X2=0 $Y2=0
cc_527 N_A1_c_714_n N_VPWR_c_756_n 0.00862f $X=8.085 $Y=1.885 $X2=0 $Y2=0
cc_528 N_A1_c_713_n N_A_722_391#_c_922_n 7.93986e-19 $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_529 N_A1_c_713_n N_A_936_391#_c_971_n 0.00902642f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_530 N_A1_c_713_n N_A_936_391#_c_974_n 0.00859469f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_531 N_A1_c_714_n N_A_936_391#_c_974_n 0.00664299f $X=8.085 $Y=1.885 $X2=0
+ $Y2=0
cc_532 N_A1_M1015_g N_VGND_c_1028_n 0.00278247f $X=7.64 $Y=0.69 $X2=0 $Y2=0
cc_533 N_A1_M1025_g N_VGND_c_1028_n 0.00278271f $X=8.1 $Y=0.69 $X2=0 $Y2=0
cc_534 N_A1_M1015_g N_VGND_c_1029_n 0.00354264f $X=7.64 $Y=0.69 $X2=0 $Y2=0
cc_535 N_A1_M1025_g N_VGND_c_1029_n 0.00357524f $X=8.1 $Y=0.69 $X2=0 $Y2=0
cc_536 N_A1_M1015_g N_A_709_119#_c_1124_n 0.0144407f $X=7.64 $Y=0.69 $X2=0 $Y2=0
cc_537 N_A1_M1025_g N_A_709_119#_c_1124_n 0.00220281f $X=8.1 $Y=0.69 $X2=0 $Y2=0
cc_538 N_A1_c_711_n N_A_709_119#_c_1124_n 0.054688f $X=8.01 $Y=1.615 $X2=0 $Y2=0
cc_539 N_A1_c_712_n N_A_709_119#_c_1124_n 0.00440863f $X=8.085 $Y=1.667 $X2=0
+ $Y2=0
cc_540 N_A1_M1015_g N_A_709_119#_c_1125_n 0.00268042f $X=7.64 $Y=0.69 $X2=0
+ $Y2=0
cc_541 N_A1_M1025_g N_A_709_119#_c_1125_n 0.00201605f $X=8.1 $Y=0.69 $X2=0 $Y2=0
cc_542 N_VPWR_M1011_d N_X_c_861_n 0.00505868f $X=1.75 $Y=1.84 $X2=0 $Y2=0
cc_543 N_VPWR_M1007_s N_A_722_391#_c_921_n 0.0120149f $X=4.06 $Y=1.955 $X2=0
+ $Y2=0
cc_544 N_VPWR_M1020_d N_A_722_391#_c_921_n 0.00917381f $X=5.13 $Y=1.955 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_760_n N_A_722_391#_c_921_n 0.0256575f $X=4.295 $Y=2.94 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_761_n N_A_722_391#_c_921_n 0.0193995f $X=5.365 $Y=2.94 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_764_n N_A_722_391#_c_921_n 0.00242035f $X=4.13 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_766_n N_A_722_391#_c_921_n 0.0088241f $X=5.2 $Y=3.33 $X2=0 $Y2=0
cc_549 N_VPWR_c_769_n N_A_722_391#_c_921_n 0.00253166f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_756_n N_A_722_391#_c_921_n 0.0298931f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_551 N_VPWR_c_769_n N_A_722_391#_c_922_n 0.0547133f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_552 N_VPWR_c_756_n N_A_722_391#_c_922_n 0.0466882f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_759_n N_A_722_391#_c_923_n 0.00758149f $X=3.225 $Y=3 $X2=0 $Y2=0
cc_554 N_VPWR_c_760_n N_A_722_391#_c_923_n 0.0132043f $X=4.295 $Y=2.94 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_764_n N_A_722_391#_c_923_n 0.0108296f $X=4.13 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_756_n N_A_722_391#_c_923_n 0.00907338f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_761_n N_A_722_391#_c_924_n 0.0156058f $X=5.365 $Y=2.94 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_769_n N_A_722_391#_c_924_n 0.00737699f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_756_n N_A_722_391#_c_924_n 0.0061588f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_560 N_VPWR_M1020_d N_A_936_391#_c_970_n 0.0142859f $X=5.13 $Y=1.955 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_756_n N_A_936_391#_c_971_n 0.020425f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_562 N_VPWR_c_769_n N_A_936_391#_c_974_n 0.0144379f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_563 N_VPWR_c_756_n N_A_936_391#_c_974_n 0.0119346f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_564 N_X_c_857_n N_VGND_c_1016_n 0.00100635f $X=1.475 $Y=1.37 $X2=0 $Y2=0
cc_565 N_X_c_858_n N_VGND_c_1016_n 0.00272557f $X=1.475 $Y=0.535 $X2=0 $Y2=0
cc_566 N_X_c_858_n N_VGND_c_1017_n 0.0270562f $X=1.475 $Y=0.535 $X2=0 $Y2=0
cc_567 N_X_c_860_n N_VGND_c_1017_n 0.0508519f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_568 N_X_c_861_n N_VGND_c_1017_n 0.0192123f $X=2.33 $Y=1.625 $X2=0 $Y2=0
cc_569 N_X_c_860_n N_VGND_c_1018_n 0.0702289f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_570 N_X_c_858_n N_VGND_c_1024_n 0.0134715f $X=1.475 $Y=0.535 $X2=0 $Y2=0
cc_571 N_X_c_860_n N_VGND_c_1026_n 0.017052f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_572 N_X_c_858_n N_VGND_c_1029_n 0.0106052f $X=1.475 $Y=0.535 $X2=0 $Y2=0
cc_573 N_X_c_860_n N_VGND_c_1029_n 0.0135629f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_574 N_A_722_391#_c_921_n N_A_936_391#_M1000_s 0.00540816f $X=5.62 $Y=2.52
+ $X2=-0.19 $Y2=1.66
cc_575 N_A_722_391#_c_922_n N_A_936_391#_c_970_n 0.00682381f $X=6.95 $Y=2.805
+ $X2=0 $Y2=0
cc_576 N_A_722_391#_c_924_n N_A_936_391#_c_970_n 0.0139328f $X=5.705 $Y=2.52
+ $X2=0 $Y2=0
cc_577 N_A_722_391#_M1004_d N_A_936_391#_c_971_n 0.00375445f $X=6.8 $Y=1.96
+ $X2=0 $Y2=0
cc_578 N_A_722_391#_c_922_n N_A_936_391#_c_971_n 0.0591194f $X=6.95 $Y=2.805
+ $X2=0 $Y2=0
cc_579 N_A_722_391#_c_921_n N_A_936_391#_c_972_n 0.0576661f $X=5.62 $Y=2.52
+ $X2=0 $Y2=0
cc_580 N_A_722_391#_c_922_n N_A_936_391#_c_973_n 0.0137316f $X=6.95 $Y=2.805
+ $X2=0 $Y2=0
cc_581 N_A_722_391#_c_924_n N_A_936_391#_c_973_n 0.0079066f $X=5.705 $Y=2.52
+ $X2=0 $Y2=0
cc_582 N_A_722_391#_c_922_n N_A_936_391#_c_974_n 0.0077481f $X=6.95 $Y=2.805
+ $X2=0 $Y2=0
cc_583 N_A_936_391#_c_972_n N_A_709_119#_c_1126_n 0.00364025f $X=5.14 $Y=2.1
+ $X2=0 $Y2=0
cc_584 N_VGND_c_1018_n N_A_709_119#_c_1122_n 0.0287269f $X=3.09 $Y=0.535 $X2=0
+ $Y2=0
cc_585 N_VGND_c_1019_n N_A_709_119#_c_1122_n 0.0075028f $X=4.02 $Y=0 $X2=0 $Y2=0
cc_586 N_VGND_c_1020_n N_A_709_119#_c_1122_n 0.0138611f $X=4.255 $Y=0.74 $X2=0
+ $Y2=0
cc_587 N_VGND_c_1029_n N_A_709_119#_c_1122_n 0.00907938f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_1018_n N_A_709_119#_c_1123_n 0.00939066f $X=3.09 $Y=0.535 $X2=0
+ $Y2=0
cc_589 N_VGND_M1010_s N_A_709_119#_c_1124_n 0.00335654f $X=5.115 $Y=0.595 $X2=0
+ $Y2=0
cc_590 N_VGND_M1024_s N_A_709_119#_c_1126_n 0.00519037f $X=4.045 $Y=0.595 $X2=0
+ $Y2=0
cc_591 N_VGND_c_1020_n N_A_709_119#_c_1126_n 0.0298247f $X=4.255 $Y=0.74 $X2=0
+ $Y2=0
cc_592 N_VGND_M1010_s N_A_709_119#_c_1127_n 0.00207907f $X=5.115 $Y=0.595 $X2=0
+ $Y2=0
cc_593 N_VGND_c_1029_n N_A_937_119#_c_1182_n 0.00702266f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_c_1020_n N_A_937_119#_c_1183_n 0.0132163f $X=4.255 $Y=0.74 $X2=0
+ $Y2=0
cc_595 N_VGND_c_1021_n N_A_937_119#_c_1183_n 7.70571e-19 $X=5.37 $Y=0.5 $X2=0
+ $Y2=0
cc_596 N_VGND_c_1027_n N_A_937_119#_c_1183_n 0.0070895f $X=5.17 $Y=0 $X2=0 $Y2=0
cc_597 N_VGND_c_1029_n N_A_937_119#_c_1183_n 0.00875466f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_M1010_s N_A_937_119#_c_1188_n 0.00778741f $X=5.115 $Y=0.595 $X2=0
+ $Y2=0
cc_599 N_VGND_c_1021_n N_A_937_119#_c_1188_n 0.0318174f $X=5.37 $Y=0.5 $X2=0
+ $Y2=0
cc_600 N_VGND_c_1027_n N_A_937_119#_c_1188_n 0.00195503f $X=5.17 $Y=0 $X2=0
+ $Y2=0
cc_601 N_VGND_c_1029_n N_A_937_119#_c_1188_n 0.005356f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_M1010_s N_A_937_119#_c_1184_n 0.00137378f $X=5.115 $Y=0.595 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1028_n N_A_937_119#_c_1184_n 0.00122935f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1029_n N_A_937_119#_c_1184_n 0.00198148f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_605 N_A_709_119#_c_1126_n N_A_937_119#_M1005_d 0.00176461f $X=5.155 $Y=1.187
+ $X2=-0.19 $Y2=-0.245
cc_606 N_A_709_119#_c_1126_n N_A_937_119#_c_1183_n 0.0161925f $X=5.155 $Y=1.187
+ $X2=0 $Y2=0
cc_607 N_A_709_119#_c_1124_n N_A_937_119#_c_1188_n 0.0115278f $X=7.77 $Y=1.195
+ $X2=0 $Y2=0
cc_608 N_A_709_119#_c_1126_n N_A_937_119#_c_1188_n 0.0196564f $X=5.155 $Y=1.187
+ $X2=0 $Y2=0
cc_609 N_A_709_119#_c_1124_n N_A_937_119#_c_1184_n 0.089963f $X=7.77 $Y=1.195
+ $X2=0 $Y2=0
cc_610 N_A_709_119#_c_1124_n N_A_937_119#_c_1199_n 0.0208323f $X=7.77 $Y=1.195
+ $X2=0 $Y2=0
