* NGSPICE file created from sky130_fd_sc_hs__or4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4_2 A B C D VGND VNB VPB VPWR X
M1000 X a_85_392# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=8.628e+11p ps=6.04e+06u
M1001 VPWR a_85_392# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_174_392# D a_85_392# VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=2.95e+11p ps=2.59e+06u
M1003 VPWR A a_342_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=4.3e+11p ps=2.86e+06u
M1004 a_258_392# C a_174_392# VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 a_85_392# B VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=1.24458e+12p ps=9.28e+06u
M1006 X a_85_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1007 a_85_392# D VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A a_85_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_85_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_85_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_342_392# B a_258_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

