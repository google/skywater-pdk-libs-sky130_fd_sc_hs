# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__clkinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.350000 5.715000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.242400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.285000 1.010000 6.115000 1.180000 ;
        RECT 0.285000 1.180000 0.455000 1.950000 ;
        RECT 0.285000 1.950000 6.115000 2.120000 ;
        RECT 0.590000 2.120000 0.920000 2.980000 ;
        RECT 0.615000 0.460000 2.625000 1.010000 ;
        RECT 1.540000 2.120000 1.870000 2.980000 ;
        RECT 2.490000 2.120000 2.820000 2.980000 ;
        RECT 3.295000 0.445000 3.625000 1.010000 ;
        RECT 3.440000 2.120000 3.770000 2.980000 ;
        RECT 4.295000 0.445000 4.625000 1.010000 ;
        RECT 4.390000 2.120000 4.720000 2.980000 ;
        RECT 5.295000 0.445000 5.625000 1.010000 ;
        RECT 5.340000 2.120000 5.670000 2.980000 ;
        RECT 5.885000 1.180000 6.115000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 6.240000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 6.430000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.775000 ;
      RECT 0.115000  2.290000 0.390000 3.245000 ;
      RECT 1.120000  2.290000 1.370000 3.245000 ;
      RECT 2.070000  2.290000 2.320000 3.245000 ;
      RECT 2.795000  0.085000 3.125000 0.775000 ;
      RECT 3.020000  2.290000 3.270000 3.245000 ;
      RECT 3.795000  0.085000 4.125000 0.775000 ;
      RECT 3.970000  2.290000 4.220000 3.245000 ;
      RECT 4.795000  0.085000 5.125000 0.775000 ;
      RECT 4.920000  2.290000 5.170000 3.245000 ;
      RECT 5.795000  0.085000 6.125000 0.775000 ;
      RECT 5.870000  2.290000 6.120000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__clkinv_8
END LIBRARY
