* NGSPICE file created from sky130_fd_sc_hs__o41a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_523_124# A4 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.1456e+12p pd=1.126e+07u as=1.69995e+12p ps=1.463e+07u
M1001 a_851_368# A3 a_762_368# VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=1.0528e+12p ps=8.6e+06u
M1002 a_762_368# A3 a_851_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_523_124# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_110_48# A4 a_851_368# VPB pshort w=1.12e+06u l=150000u
+  ad=5.992e+11p pd=5.14e+06u as=0p ps=0u
M1005 a_523_124# B1 a_110_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 a_1213_368# A2 a_762_368# VPB pshort w=1.12e+06u l=150000u
+  ad=7.28e+11p pd=5.78e+06u as=0p ps=0u
M1007 VPWR A1 a_1213_368# VPB pshort w=1.12e+06u l=150000u
+  ad=1.6953e+12p pd=1.387e+07u as=0p ps=0u
M1008 a_523_124# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_110_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1010 a_523_124# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A1 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_110_48# B1 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_110_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A3 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_110_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_110_48# B1 VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A2 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_762_368# A2 a_1213_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_110_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1020 VPWR B1 a_110_48# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1213_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_110_48# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_110_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_110_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_110_48# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_851_368# A4 a_110_48# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A4 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

