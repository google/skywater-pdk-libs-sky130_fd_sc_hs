* NGSPICE file created from sky130_fd_sc_hs__a311oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=7.178e+11p ps=4.9e+06u
M1001 a_127_368# A3 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=1.344e+12p pd=1.136e+07u as=1.3216e+12p ps=1.132e+07u
M1002 VPWR A3 a_127_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_127_368# A2 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_127_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_127_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_45_74# A2 a_300_74# VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=4.144e+11p ps=4.08e+06u
M1007 VPWR A1 a_127_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_45_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A3 a_45_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_127_368# B1 a_692_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=9.52e+11p ps=8.42e+06u
M1011 Y A1 a_300_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_692_368# B1 a_127_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C1 a_692_368# VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1014 a_300_74# A2 a_45_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_692_368# C1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_300_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

