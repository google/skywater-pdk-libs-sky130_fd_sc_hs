* File: sky130_fd_sc_hs__sdfrtp_1.pex.spice
* Created: Thu Aug 27 21:08:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%SCE 2 5 7 9 11 12 14 17 19 22 23 27 28 29
+ 37 43 52 54
c87 37 0 9.7872e-20 $X=0.96 $Y=1.67
c88 22 0 2.01624e-19 $X=2.56 $Y=1.425
r89 43 52 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=1.623 $Y=1.662
+ $X2=1.68 $Y2=1.662
r90 37 39 6.6128 $w=3.28e-07 $l=4.5e-08 $layer=POLY_cond $X=0.96 $Y=1.67
+ $X2=1.005 $Y2=1.67
r91 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.96
+ $Y=1.67 $X2=0.96 $Y2=1.67
r92 35 37 66.8628 $w=3.28e-07 $l=4.55e-07 $layer=POLY_cond $X=0.505 $Y=1.67
+ $X2=0.96 $Y2=1.67
r93 34 35 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.67
+ $X2=0.505 $Y2=1.67
r94 29 54 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.795 $Y2=1.662
r95 29 52 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.68 $Y2=1.662
r96 29 43 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.623 $Y2=1.662
r97 28 29 13.6623 $w=3.43e-07 $l=4.09e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=1.609 $Y2=1.662
r98 28 38 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=0.96 $Y2=1.662
r99 27 38 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=1.662
+ $X2=0.96 $Y2=1.662
r100 23 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.56 $Y=1.425
+ $X2=2.56 $Y2=1.26
r101 22 25 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.56 $Y=1.425
+ $X2=2.56 $Y2=1.575
r102 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.425 $X2=2.56 $Y2=1.425
r103 19 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=1.575
+ $X2=2.56 $Y2=1.575
r104 19 54 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.395 $Y=1.575
+ $X2=1.795 $Y2=1.575
r105 17 41 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.65 $Y=0.615
+ $X2=2.65 $Y2=1.26
r106 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.005 $Y=2.245
+ $X2=1.005 $Y2=2.64
r107 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.005 $Y=2.155
+ $X2=1.005 $Y2=2.245
r108 10 39 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.835
+ $X2=1.005 $Y2=1.67
r109 10 11 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=1.835
+ $X2=1.005 $Y2=2.155
r110 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r111 3 34 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=1.67
r112 3 5 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=0.65
r113 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.155
+ $X2=0.505 $Y2=2.245
r114 1 35 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=1.67
r115 1 2 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_27_88# 1 2 7 9 12 14 17 20 23 25 29 31 32
+ 34 35 37 38 42
c84 37 0 9.7872e-20 $X=1.21 $Y=1.1
c85 7 0 3.56444e-20 $X=1.485 $Y=0.935
r86 37 40 1.99058 $w=3.28e-07 $l=5.7e-08 $layer=LI1_cond $X=1.21 $Y=1.1 $X2=1.21
+ $Y2=1.157
r87 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.1 $X2=1.21 $Y2=1.1
r88 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.54
+ $Y=1.995 $X2=2.54 $Y2=1.995
r89 29 42 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=2.207 $Y=2.002
+ $X2=2.035 $Y2=2.002
r90 29 31 11.1236 $w=3.43e-07 $l=3.33e-07 $layer=LI1_cond $X=2.207 $Y=2.002
+ $X2=2.54 $Y2=2.002
r91 28 35 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=0.28 $Y2=2.09
r92 28 42 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=2.035 $Y2=2.09
r93 26 34 1.25797 $w=2.15e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.157
+ $X2=0.24 $Y2=1.157
r94 25 40 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=1.157
+ $X2=1.21 $Y2=1.157
r95 25 26 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=1.157
+ $X2=0.365 $Y2=1.157
r96 21 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.09
r97 21 23 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.465
r98 20 35 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.005
+ $X2=0.28 $Y2=2.09
r99 19 34 5.26796 $w=2.1e-07 $l=1.26428e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.24 $Y2=1.157
r100 19 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.2 $Y2=2.005
r101 15 34 5.26796 $w=2.1e-07 $l=1.07e-07 $layer=LI1_cond $X=0.24 $Y=1.05
+ $X2=0.24 $Y2=1.157
r102 15 17 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=1.05 $X2=0.24
+ $Y2=0.65
r103 12 32 19.685 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.615 $Y=2.245
+ $X2=2.615 $Y2=2.037
r104 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.615 $Y=2.245
+ $X2=2.615 $Y2=2.64
r105 7 38 50.0189 $w=2.65e-07 $l=3.47851e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.21 $Y2=1.1
r106 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.615
r107 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r108 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.44 $X2=0.28 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%D 1 3 5 7 10 11 15 17 20 21 22
c54 15 0 5.92372e-20 $X=1.845 $Y=1.515
c55 5 0 1.42386e-19 $X=1.69 $Y=2.075
r56 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.1
+ $X2=1.935 $Y2=1.265
r57 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.1
+ $X2=1.935 $Y2=0.935
r58 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.1 $X2=1.935 $Y2=1.1
r59 17 21 6.7033 $w=4.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.037
+ $X2=1.935 $Y2=1.037
r60 13 15 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.845 $Y2=1.515
r61 11 12 80.8418 $w=1.58e-07 $l=2.65e-07 $layer=POLY_cond $X=1.425 $Y=2.16
+ $X2=1.69 $Y2=2.16
r62 10 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.875 $Y=0.615
+ $X2=1.875 $Y2=0.935
r63 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.44
+ $X2=1.845 $Y2=1.515
r64 7 23 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.845 $Y=1.44
+ $X2=1.845 $Y2=1.265
r65 5 12 4.07462 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.69 $Y=2.075
+ $X2=1.69 $Y2=2.16
r66 4 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.59 $X2=1.69
+ $Y2=1.515
r67 4 5 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.69 $Y=1.59 $X2=1.69
+ $Y2=2.075
r68 1 11 4.07462 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.425 $Y=2.245
+ $X2=1.425 $Y2=2.16
r69 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.425 $Y=2.245
+ $X2=1.425 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%SCD 1 3 6 10 11 12 16
c44 6 0 3.56444e-20 $X=3.04 $Y=0.615
r45 11 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.035
r46 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.11
+ $Y=1.605 $X2=3.11 $Y2=1.605
r47 10 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.11 $Y=1.945
+ $X2=3.11 $Y2=1.605
r48 9 16 43.0552 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.44
+ $X2=3.11 $Y2=1.605
r49 6 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.04 $Y=0.615
+ $X2=3.04 $Y2=1.44
r50 1 10 55.1908 $w=2.62e-07 $l=3.3541e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.11 $Y2=1.945
r51 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.035 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%RESET_B 1 3 6 8 10 11 12 14 15 17 20 23 25
+ 26 28 33 35 36 37 38 45 46 49 50 53 61 62
c212 37 0 1.37312e-19 $X=10.655 $Y=2.035
c213 33 0 6.31244e-20 $X=10.715 $Y=1.375
c214 20 0 5.21422e-20 $X=10.6 $Y=0.58
c215 12 0 8.22544e-20 $X=7.375 $Y=1.16
c216 8 0 1.64601e-19 $X=7.3 $Y=1.085
c217 6 0 8.6114e-20 $X=3.655 $Y=0.615
r218 60 62 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=10.805 $Y=1.985
+ $X2=10.885 $Y2=1.985
r219 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.805
+ $Y=1.985 $X2=10.805 $Y2=1.985
r220 57 60 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.715 $Y=1.985
+ $X2=10.805 $Y2=1.985
r221 53 55 42.6489 $w=3.56e-07 $l=3.15e-07 $layer=POLY_cond $X=7.685 $Y=2.022
+ $X2=8 $Y2=2.022
r222 52 53 2.0309 $w=3.56e-07 $l=1.5e-08 $layer=POLY_cond $X=7.67 $Y=2.022
+ $X2=7.685 $Y2=2.022
r223 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r224 46 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r225 45 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8 $Y=1.98
+ $X2=8 $Y2=1.98
r226 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r227 40 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r228 38 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r229 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r230 37 38 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r231 36 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r232 35 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r233 35 36 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r234 31 33 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=10.6 $Y=1.375
+ $X2=10.715 $Y2=1.375
r235 30 49 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.73 $Y=1.995
+ $X2=3.95 $Y2=1.995
r236 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.885 $Y=2.465
+ $X2=10.885 $Y2=2.75
r237 25 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.885 $Y=2.375
+ $X2=10.885 $Y2=2.465
r238 24 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.885 $Y=2.15
+ $X2=10.885 $Y2=1.985
r239 24 25 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=10.885 $Y=2.15
+ $X2=10.885 $Y2=2.375
r240 23 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.715 $Y=1.82
+ $X2=10.715 $Y2=1.985
r241 22 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.715 $Y=1.45
+ $X2=10.715 $Y2=1.375
r242 22 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.715 $Y=1.45
+ $X2=10.715 $Y2=1.82
r243 18 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.6 $Y2=1.375
r244 18 20 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.6 $Y2=0.58
r245 15 53 23.0368 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.685 $Y=2.23
+ $X2=7.685 $Y2=2.022
r246 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.685 $Y=2.23
+ $X2=7.685 $Y2=2.515
r247 14 52 23.0368 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.67 $Y=1.815
+ $X2=7.67 $Y2=2.022
r248 13 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.67 $Y=1.235
+ $X2=7.67 $Y2=1.815
r249 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.595 $Y=1.16
+ $X2=7.67 $Y2=1.235
r250 11 12 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=7.595 $Y=1.16
+ $X2=7.375 $Y2=1.16
r251 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.3 $Y=1.085
+ $X2=7.375 $Y2=1.16
r252 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.3 $Y=1.085 $X2=7.3
+ $Y2=0.8
r253 4 30 45.8367 $w=1.79e-07 $l=1.80748e-07 $layer=POLY_cond $X=3.655 $Y=1.83
+ $X2=3.622 $Y2=1.995
r254 4 6 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.655 $Y=1.83
+ $X2=3.655 $Y2=0.615
r255 1 30 68.725 $w=1.79e-07 $l=2.5836e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.622 $Y2=1.995
r256 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%CLK 1 3 6 9 12 15 22
c52 6 0 2.38973e-19 $X=4.665 $Y=0.74
r53 15 22 3.70473 $w=4.08e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.385
+ $X2=4.195 $Y2=1.385
r54 12 22 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.475 $Y=1.425
+ $X2=4.195 $Y2=1.425
r55 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.475
+ $Y=1.425 $X2=4.475 $Y2=1.425
r56 9 13 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=4.555 $Y=1.425
+ $X2=4.475 $Y2=1.425
r57 4 9 45.1689 $w=1.83e-07 $l=1.73767e-07 $layer=POLY_cond $X=4.665 $Y=1.26
+ $X2=4.647 $Y2=1.425
r58 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=4.665 $Y=1.26
+ $X2=4.665 $Y2=0.74
r59 1 9 91.2618 $w=1.83e-07 $l=3.40999e-07 $layer=POLY_cond $X=4.645 $Y=1.765
+ $X2=4.647 $Y2=1.425
r60 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_1034_368# 1 2 8 9 11 12 16 18 20 22 23 25
+ 29 31 32 33 34 36 40 41 42 44 45 46 48 50 51 53 56 64 65 67 72
c213 67 0 1.29298e-19 $X=6.065 $Y=1.65
c214 65 0 1.39473e-19 $X=9.33 $Y=1.105
c215 56 0 1.36239e-19 $X=5.385 $Y=1.13
c216 42 0 1.07934e-19 $X=7.22 $Y=0.665
c217 33 0 1.02734e-19 $X=5.62 $Y=0.34
c218 16 0 6.15336e-20 $X=6.52 $Y=0.8
c219 9 0 1.93993e-19 $X=6.135 $Y=2.21
r220 64 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.105
+ $X2=9.085 $Y2=1.105
r221 63 65 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.25 $Y=1.105 $X2=9.33
+ $Y2=1.105
r222 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.25
+ $Y=1.105 $X2=9.25 $Y2=1.105
r223 60 63 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=9.15 $Y=1.105
+ $X2=9.25 $Y2=1.105
r224 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.81
+ $Y=2.215 $X2=9.81 $Y2=2.215
r225 51 53 17.8516 $w=2.53e-07 $l=3.95e-07 $layer=LI1_cond $X=9.415 $Y=2.252
+ $X2=9.81 $Y2=2.252
r226 50 51 7.17723 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=9.33 $Y=2.125
+ $X2=9.415 $Y2=2.252
r227 49 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.33 $Y=1.27
+ $X2=9.33 $Y2=1.105
r228 49 50 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=9.33 $Y=1.27
+ $X2=9.33 $Y2=2.125
r229 48 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=0.94
+ $X2=9.15 $Y2=1.105
r230 47 48 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=9.15 $Y=0.425
+ $X2=9.15 $Y2=0.94
r231 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.065 $Y=0.34
+ $X2=9.15 $Y2=0.425
r232 45 46 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=9.065 $Y=0.34
+ $X2=8.1 $Y2=0.34
r233 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.1 $Y2=0.34
r234 43 44 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.015 $Y2=0.58
r235 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=8.015 $Y2=0.58
r236 41 42 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=7.22 $Y2=0.665
r237 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.135 $Y=0.58
+ $X2=7.22 $Y2=0.665
r238 39 40 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.135 $Y=0.425
+ $X2=7.135 $Y2=0.58
r239 37 70 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=1.71
+ $X2=6.065 $Y2=1.875
r240 37 67 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.065 $Y=1.71
+ $X2=6.065 $Y2=1.65
r241 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.71 $X2=6.065 $Y2=1.71
r242 34 59 10.9942 $w=3.44e-07 $l=4.1028e-07 $layer=LI1_cond $X=5.62 $Y=1.71
+ $X2=5.387 $Y2=2.02
r243 34 36 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.62 $Y=1.71
+ $X2=6.065 $Y2=1.71
r244 32 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=7.135 $Y2=0.425
r245 32 33 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=5.62 $Y2=0.34
r246 31 34 8.97475 $w=3.44e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.535 $Y=1.545
+ $X2=5.62 $Y2=1.71
r247 31 56 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.535 $Y=1.545
+ $X2=5.535 $Y2=1.13
r248 27 56 11.119 $w=4.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.385 $Y=0.895
+ $X2=5.385 $Y2=1.13
r249 27 29 9.67042 $w=4.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.385 $Y=0.895
+ $X2=5.385 $Y2=0.515
r250 26 33 8.97637 $w=1.7e-07 $l=2.74226e-07 $layer=LI1_cond $X=5.385 $Y=0.425
+ $X2=5.62 $Y2=0.34
r251 26 29 2.29036 $w=4.68e-07 $l=9e-08 $layer=LI1_cond $X=5.385 $Y=0.425
+ $X2=5.385 $Y2=0.515
r252 23 54 52.063 $w=3.03e-07 $l=2.86356e-07 $layer=POLY_cond $X=9.89 $Y=2.465
+ $X2=9.812 $Y2=2.215
r253 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.89 $Y=2.465
+ $X2=9.89 $Y2=2.75
r254 22 72 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=8.725 $Y=1.16
+ $X2=9.085 $Y2=1.16
r255 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.725 $Y2=1.16
r256 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.65 $Y2=0.69
r257 14 16 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=6.52 $Y=1.575
+ $X2=6.52 $Y2=0.8
r258 13 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.65
+ $X2=6.065 $Y2=1.65
r259 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.445 $Y=1.65
+ $X2=6.52 $Y2=1.575
r260 12 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.445 $Y=1.65
+ $X2=6.23 $Y2=1.65
r261 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.135 $Y=2.21
+ $X2=6.135 $Y2=2.495
r262 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.135 $Y=2.12 $X2=6.135
+ $Y2=2.21
r263 8 70 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=6.135 $Y=2.12
+ $X2=6.135 $Y2=1.875
r264 2 59 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.84 $X2=5.32 $Y2=2.02
r265 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.175
+ $Y=0.37 $X2=5.315 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_1367_92# 1 2 9 12 13 15 18 19 21 22 25 27
+ 32 34
c109 22 0 8.22544e-20 $X=7.325 $Y=1.005
c110 9 0 1.57288e-19 $X=6.91 $Y=0.8
r111 35 37 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=6.91 $Y=1.64
+ $X2=7.06 $Y2=1.64
r112 27 29 29.2227 $w=2.78e-07 $l=7.1e-07 $layer=LI1_cond $X=8.865 $Y=1.88
+ $X2=8.865 $Y2=2.59
r113 25 34 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=8.865 $Y=1.855
+ $X2=8.865 $Y2=1.715
r114 25 27 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=8.865 $Y=1.855
+ $X2=8.865 $Y2=1.88
r115 23 32 12.3649 $w=3.7e-07 $l=4.83348e-07 $layer=LI1_cond $X=8.81 $Y=1.09
+ $X2=8.435 $Y2=0.842
r116 23 34 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=8.81 $Y=1.09
+ $X2=8.81 $Y2=1.715
r117 21 32 9.03936 $w=3.7e-07 $l=2.32637e-07 $layer=LI1_cond $X=8.27 $Y=1.005
+ $X2=8.435 $Y2=0.842
r118 21 22 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=8.27 $Y=1.005
+ $X2=7.325 $Y2=1.005
r119 19 37 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=7.185 $Y=1.64
+ $X2=7.06 $Y2=1.64
r120 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.185
+ $Y=1.64 $X2=7.185 $Y2=1.64
r121 16 22 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=7.187 $Y=1.09
+ $X2=7.325 $Y2=1.005
r122 16 18 23.0489 $w=2.73e-07 $l=5.5e-07 $layer=LI1_cond $X=7.187 $Y=1.09
+ $X2=7.187 $Y2=1.64
r123 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.06 $Y=2.23
+ $X2=7.06 $Y2=2.515
r124 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.06 $Y=2.14 $X2=7.06
+ $Y2=2.23
r125 11 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.06 $Y=1.805
+ $X2=7.06 $Y2=1.64
r126 11 12 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=7.06 $Y=1.805
+ $X2=7.06 $Y2=2.14
r127 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=1.64
r128 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=0.8
r129 2 29 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.735 $X2=8.92 $Y2=2.59
r130 2 27 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.735 $X2=8.92 $Y2=1.88
r131 1 32 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.37 $X2=8.435 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_1233_118# 1 2 3 12 14 16 18 19 23 26 27
+ 30 31 33 34 37 41
c134 41 0 1.93993e-19 $X=6.795 $Y=2.522
c135 30 0 7.00504e-20 $X=7.58 $Y=2.32
c136 26 0 3.48885e-19 $X=6.795 $Y=2.32
c137 23 0 1.49497e-20 $X=6.71 $Y=0.945
r138 37 39 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.305 $Y=0.81
+ $X2=6.305 $Y2=0.945
r139 34 46 16.6207 $w=3.19e-07 $l=1.1e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.52
r140 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.15
+ $Y=1.41 $X2=8.15 $Y2=1.41
r141 31 33 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=7.665 $Y=1.417
+ $X2=8.15 $Y2=1.417
r142 30 44 12.781 $w=3.15e-07 $l=4.22918e-07 $layer=LI1_cond $X=7.58 $Y=2.32
+ $X2=7.91 $Y2=2.532
r143 29 31 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.665 $Y2=1.417
r144 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.58 $Y2=2.32
r145 28 41 3.64284 $w=2.55e-07 $l=1.53734e-07 $layer=LI1_cond $X=6.88 $Y=2.405
+ $X2=6.795 $Y2=2.522
r146 27 30 5.86024 $w=3.15e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=7.58 $Y2=2.32
r147 27 28 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=6.88 $Y2=2.405
r148 26 41 2.83584 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=6.795 $Y=2.32
+ $X2=6.795 $Y2=2.522
r149 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=6.795 $Y=1.03
+ $X2=6.795 $Y2=2.32
r150 24 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.47 $Y=0.945
+ $X2=6.305 $Y2=0.945
r151 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.71 $Y=0.945
+ $X2=6.795 $Y2=1.03
r152 23 24 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.71 $Y=0.945
+ $X2=6.47 $Y2=0.945
r153 19 41 3.64284 $w=2.55e-07 $l=1.0015e-07 $layer=LI1_cond $X=6.71 $Y=2.555
+ $X2=6.795 $Y2=2.522
r154 19 21 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=6.71 $Y=2.555
+ $X2=6.415 $Y2=2.555
r155 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.695 $Y=1.66
+ $X2=8.695 $Y2=2.235
r156 15 46 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.315 $Y=1.52
+ $X2=8.15 $Y2=1.52
r157 14 16 26.9307 $w=1.5e-07 $l=1.79444e-07 $layer=POLY_cond $X=8.605 $Y=1.52
+ $X2=8.695 $Y2=1.66
r158 14 15 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.605 $Y=1.52
+ $X2=8.315 $Y2=1.52
r159 10 34 38.5462 $w=3.19e-07 $l=1.96914e-07 $layer=POLY_cond $X=8.22 $Y=1.245
+ $X2=8.15 $Y2=1.41
r160 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.22 $Y=1.245
+ $X2=8.22 $Y2=0.69
r161 3 44 600 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.305 $X2=7.91 $Y2=2.53
r162 2 21 600 $w=1.7e-07 $l=3.5812e-07 $layer=licon1_PDIFF $count=1 $X=6.21
+ $Y=2.285 $X2=6.415 $Y2=2.555
r163 1 37 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=6.165
+ $Y=0.59 $X2=6.305 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_855_368# 1 2 7 9 10 12 13 16 17 19 20 23
+ 25 26 27 29 30 32 33 37 38 39 41 44 46 47 50 54 56 57 58 61 63 64 72
c202 44 0 2.96321e-20 $X=9.785 $Y=0.58
c203 38 0 1.09841e-19 $X=9.625 $Y=1.585
c204 23 0 1.49497e-20 $X=6.09 $Y=0.8
c205 7 0 6.15093e-20 $X=5.095 $Y=1.765
r206 73 75 33.4949 $w=2.95e-07 $l=2.05e-07 $layer=POLY_cond $X=5.115 $Y=1.465
+ $X2=5.115 $Y2=1.26
r207 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.465 $X2=5.115 $Y2=1.465
r208 69 72 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.895 $Y=1.465
+ $X2=5.115 $Y2=1.465
r209 64 67 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.46 $Y=1.905
+ $X2=4.46 $Y2=2.02
r210 62 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=1.63
+ $X2=4.895 $Y2=1.465
r211 62 63 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.895 $Y=1.63
+ $X2=4.895 $Y2=1.82
r212 61 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=1.3
+ $X2=4.895 $Y2=1.465
r213 60 61 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.895 $Y=1.09
+ $X2=4.895 $Y2=1.3
r214 59 64 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=1.905
+ $X2=4.46 $Y2=1.905
r215 58 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.81 $Y=1.905
+ $X2=4.895 $Y2=1.82
r216 58 59 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.81 $Y=1.905
+ $X2=4.585 $Y2=1.905
r217 56 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.81 $Y=1.005
+ $X2=4.895 $Y2=1.09
r218 56 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.81 $Y=1.005
+ $X2=4.535 $Y2=1.005
r219 52 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.45 $Y=0.92
+ $X2=4.535 $Y2=1.005
r220 52 54 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.45 $Y=0.92
+ $X2=4.45 $Y2=0.515
r221 48 50 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=9.7 $Y=1.045
+ $X2=9.785 $Y2=1.045
r222 42 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.785 $Y=0.97
+ $X2=9.785 $Y2=1.045
r223 42 44 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=9.785 $Y=0.97
+ $X2=9.785 $Y2=0.58
r224 40 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.7 $Y=1.12 $X2=9.7
+ $Y2=1.045
r225 40 41 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=9.7 $Y=1.12 $X2=9.7
+ $Y2=1.51
r226 38 41 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.7 $Y2=1.51
r227 38 39 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.22 $Y2=1.585
r228 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.145 $Y=2.81
+ $X2=9.145 $Y2=2.235
r229 34 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.145 $Y=1.66
+ $X2=9.22 $Y2=1.585
r230 34 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.145 $Y=1.66
+ $X2=9.145 $Y2=2.235
r231 32 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.145 $Y=2.9
+ $X2=9.145 $Y2=2.81
r232 32 33 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=9.145 $Y=2.9
+ $X2=9.145 $Y2=3.075
r233 31 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.73 $Y=3.15 $X2=6.64
+ $Y2=3.15
r234 30 33 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.055 $Y=3.15
+ $X2=9.145 $Y2=3.075
r235 30 31 1192.18 $w=1.5e-07 $l=2.325e-06 $layer=POLY_cond $X=9.055 $Y=3.15
+ $X2=6.73 $Y2=3.15
r236 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.64 $Y=2.8 $X2=6.64
+ $Y2=2.515
r237 26 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.64 $Y=3.075
+ $X2=6.64 $Y2=3.15
r238 25 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.64 $Y=2.89 $X2=6.64
+ $Y2=2.8
r239 25 26 71.9113 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=6.64 $Y=2.89
+ $X2=6.64 $Y2=3.075
r240 21 23 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=6.09 $Y=1.185
+ $X2=6.09 $Y2=0.8
r241 19 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.55 $Y=3.15 $X2=6.64
+ $Y2=3.15
r242 19 20 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.55 $Y=3.15
+ $X2=5.69 $Y2=3.15
r243 18 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.69 $Y=1.26
+ $X2=5.615 $Y2=1.26
r244 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.015 $Y=1.26
+ $X2=6.09 $Y2=1.185
r245 17 18 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=6.015 $Y=1.26
+ $X2=5.69 $Y2=1.26
r246 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=3.075
+ $X2=5.69 $Y2=3.15
r247 15 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.615 $Y=1.335
+ $X2=5.615 $Y2=1.26
r248 15 16 892.213 $w=1.5e-07 $l=1.74e-06 $layer=POLY_cond $X=5.615 $Y=1.335
+ $X2=5.615 $Y2=3.075
r249 14 75 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.28 $Y=1.26
+ $X2=5.115 $Y2=1.26
r250 13 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.54 $Y=1.26
+ $X2=5.615 $Y2=1.26
r251 13 14 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.54 $Y=1.26
+ $X2=5.28 $Y2=1.26
r252 10 75 23.8729 $w=2.95e-07 $l=8.21584e-08 $layer=POLY_cond $X=5.1 $Y=1.185
+ $X2=5.115 $Y2=1.26
r253 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.1 $Y=1.185
+ $X2=5.1 $Y2=0.74
r254 7 73 60.6356 $w=2.95e-07 $l=3.09839e-07 $layer=POLY_cond $X=5.095 $Y=1.765
+ $X2=5.115 $Y2=1.465
r255 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.095 $Y=1.765
+ $X2=5.095 $Y2=2.4
r256 2 67 600 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.84 $X2=4.42 $Y2=2.02
r257 1 54 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.305
+ $Y=0.37 $X2=4.45 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_1997_272# 1 2 9 11 12 13 15 16 20 24 26
+ 27 29 34 36 37 39
c117 34 0 6.31244e-20 $X=10.315 $Y=1.525
c118 29 0 1.53844e-19 $X=11.65 $Y=1.445
c119 16 0 6.72618e-20 $X=11.14 $Y=1.53
r120 36 37 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=11.127 $Y=2.75
+ $X2=11.127 $Y2=2.52
r121 31 34 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=10.15 $Y=1.525
+ $X2=10.315 $Y2=1.525
r122 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.15
+ $Y=1.525 $X2=10.15 $Y2=1.525
r123 28 29 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.65 $Y=0.925
+ $X2=11.65 $Y2=1.445
r124 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.65 $Y2=0.925
r125 26 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.34 $Y2=0.84
r126 25 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.31 $Y=1.53
+ $X2=11.225 $Y2=1.53
r127 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.565 $Y=1.53
+ $X2=11.65 $Y2=1.445
r128 24 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.565 $Y=1.53
+ $X2=11.31 $Y2=1.53
r129 22 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.225 $Y=1.615
+ $X2=11.225 $Y2=1.53
r130 22 37 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=11.225 $Y=1.615
+ $X2=11.225 $Y2=2.52
r131 18 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.175 $Y=0.755
+ $X2=11.34 $Y2=0.84
r132 18 20 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=11.175 $Y=0.755
+ $X2=11.175 $Y2=0.58
r133 16 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.14 $Y=1.53
+ $X2=11.225 $Y2=1.53
r134 16 34 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=11.14 $Y=1.53
+ $X2=10.315 $Y2=1.53
r135 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.31 $Y=2.465
+ $X2=10.31 $Y2=2.75
r136 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.31 $Y=2.375
+ $X2=10.31 $Y2=2.465
r137 11 32 58.2622 $w=3e-07 $l=3.69317e-07 $layer=POLY_cond $X=10.31 $Y=1.84
+ $X2=10.192 $Y2=1.525
r138 11 12 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=10.31 $Y=1.84
+ $X2=10.31 $Y2=2.375
r139 7 32 38.5519 $w=3e-07 $l=1.87029e-07 $layer=POLY_cond $X=10.145 $Y=1.36
+ $X2=10.192 $Y2=1.525
r140 7 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=10.145 $Y=1.36
+ $X2=10.145 $Y2=0.58
r141 2 36 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=2.54 $X2=11.11 $Y2=2.75
r142 1 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.37 $X2=11.175 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_1745_74# 1 2 9 12 14 15 17 18 19 20 22 24
+ 27 29 30 35 37 40 41 43 45 48 50 52
c167 50 0 5.21422e-20 $X=11.23 $Y=1.185
c168 43 0 1.05093e-19 $X=10.23 $Y=2.55
c169 12 0 1.53844e-19 $X=11.32 $Y=1.84
r170 51 56 13.6415 $w=3.18e-07 $l=9e-08 $layer=POLY_cond $X=11.23 $Y=1.145
+ $X2=11.32 $Y2=1.145
r171 50 52 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=11.23 $Y=1.185
+ $X2=11.065 $Y2=1.185
r172 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.23
+ $Y=1.185 $X2=11.23 $Y2=1.185
r173 45 47 9.9702 $w=3.48e-07 $l=2.1e-07 $layer=LI1_cond $X=9.58 $Y=0.56
+ $X2=9.58 $Y2=0.77
r174 42 43 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=10.23 $Y=1.955
+ $X2=10.23 $Y2=2.55
r175 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.145 $Y=1.87
+ $X2=10.23 $Y2=1.955
r176 40 41 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.145 $Y=1.87
+ $X2=9.755 $Y2=1.87
r177 39 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.755 $Y=1.18
+ $X2=9.67 $Y2=1.18
r178 39 52 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=9.755 $Y=1.18
+ $X2=11.065 $Y2=1.18
r179 37 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.67 $Y=1.785
+ $X2=9.755 $Y2=1.87
r180 36 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=1.265
+ $X2=9.67 $Y2=1.18
r181 36 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.67 $Y=1.265
+ $X2=9.67 $Y2=1.785
r182 35 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=1.095
+ $X2=9.67 $Y2=1.18
r183 35 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.67 $Y=1.095
+ $X2=9.67 $Y2=0.77
r184 30 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.145 $Y=2.715
+ $X2=10.23 $Y2=2.55
r185 30 32 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=10.145 $Y=2.715
+ $X2=9.56 $Y2=2.715
r186 25 27 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=11.955 $Y=1.2
+ $X2=11.955 $Y2=0.645
r187 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.92 $Y=2.045
+ $X2=11.92 $Y2=2.54
r188 21 29 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.425 $Y=1.915
+ $X2=11.335 $Y2=1.915
r189 20 22 26.9307 $w=1.5e-07 $l=1.69115e-07 $layer=POLY_cond $X=11.83 $Y=1.915
+ $X2=11.92 $Y2=2.045
r190 20 21 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=11.83 $Y=1.915
+ $X2=11.425 $Y2=1.915
r191 19 56 24.9017 $w=3.18e-07 $l=1.63248e-07 $layer=POLY_cond $X=11.395
+ $Y=1.275 $X2=11.32 $Y2=1.145
r192 18 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.88 $Y=1.275
+ $X2=11.955 $Y2=1.2
r193 18 19 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.88 $Y=1.275
+ $X2=11.395 $Y2=1.275
r194 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.335 $Y=2.465
+ $X2=11.335 $Y2=2.75
r195 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.335 $Y=2.375
+ $X2=11.335 $Y2=2.465
r196 13 29 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.335 $Y=1.99
+ $X2=11.335 $Y2=1.915
r197 13 14 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=11.335 $Y=1.99
+ $X2=11.335 $Y2=2.375
r198 12 29 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.32 $Y=1.84
+ $X2=11.335 $Y2=1.915
r199 11 56 20.3436 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=11.32 $Y=1.35
+ $X2=11.32 $Y2=1.145
r200 11 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=11.32 $Y=1.35
+ $X2=11.32 $Y2=1.84
r201 7 51 40.9245 $w=3.18e-07 $l=3.5812e-07 $layer=POLY_cond $X=10.96 $Y=0.94
+ $X2=11.23 $Y2=1.145
r202 7 9 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=10.96 $Y=0.94
+ $X2=10.96 $Y2=0.58
r203 2 32 600 $w=1.7e-07 $l=1.13737e-06 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.735 $X2=9.56 $Y2=2.715
r204 1 45 182 $w=1.7e-07 $l=9.35187e-07 $layer=licon1_NDIFF $count=1 $X=8.725
+ $Y=0.37 $X2=9.57 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_2399_424# 1 2 7 9 12 15 19 23 29 32 33
r47 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.745
+ $Y=1.465 $X2=12.745 $Y2=1.465
r48 27 33 0.189605 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=12.335 $Y=1.465
+ $X2=12.21 $Y2=1.465
r49 27 29 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=12.335 $Y=1.465
+ $X2=12.745 $Y2=1.465
r50 25 33 6.72893 $w=2.37e-07 $l=1.71377e-07 $layer=LI1_cond $X=12.197 $Y=1.63
+ $X2=12.21 $Y2=1.465
r51 25 32 24.0733 $w=2.23e-07 $l=4.7e-07 $layer=LI1_cond $X=12.197 $Y=1.63
+ $X2=12.197 $Y2=2.1
r52 21 33 6.72893 $w=2.37e-07 $l=1.65e-07 $layer=LI1_cond $X=12.21 $Y=1.3
+ $X2=12.21 $Y2=1.465
r53 21 23 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=12.21 $Y=1.3
+ $X2=12.21 $Y2=0.645
r54 19 32 6.93655 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.145 $Y=2.265
+ $X2=12.145 $Y2=2.1
r55 15 30 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=12.84 $Y=1.465
+ $X2=12.745 $Y2=1.465
r56 15 16 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.93 $Y=1.465
+ $X2=12.93 $Y2=1.3
r57 12 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.945 $Y=0.74
+ $X2=12.945 $Y2=1.3
r58 7 15 118.763 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=12.93 $Y=1.765
+ $X2=12.93 $Y2=1.465
r59 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.93 $Y=1.765
+ $X2=12.93 $Y2=2.4
r60 2 19 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=11.995
+ $Y=2.12 $X2=12.145 $Y2=2.265
r61 1 23 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=12.03
+ $Y=0.37 $X2=12.17 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 41 45 51
+ 55 61 66 67 69 70 72 73 74 76 81 93 110 116 117 120 123 126 129 132
c162 2 0 1.19423e-19 $X=3.11 $Y=2.32
r163 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r164 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r165 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r166 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r167 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r168 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r169 117 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r170 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r171 114 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.87 $Y=3.33
+ $X2=12.705 $Y2=3.33
r172 114 116 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=12.87 $Y=3.33
+ $X2=13.2 $Y2=3.33
r173 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r174 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r175 110 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.705 $Y2=3.33
r176 110 112 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.24 $Y2=3.33
r177 109 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r178 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r179 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r180 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r181 103 106 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r182 103 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r183 102 105 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r184 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r185 100 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.47 $Y2=3.33
r186 100 102 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.88 $Y2=3.33
r187 99 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r188 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r189 95 98 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r190 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r191 93 126 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=7.372 $Y2=3.33
r192 93 98 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=6.96 $Y2=3.33
r193 92 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r194 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r195 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r196 89 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r197 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r198 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r199 86 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r200 86 88 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r201 85 124 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r202 85 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r203 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r204 82 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r205 82 84 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r206 81 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r207 81 84 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.2 $Y2=3.33
r208 79 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r209 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r210 76 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r211 76 78 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r212 74 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r213 74 96 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=5.04 $Y2=3.33
r214 72 108 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=11.48 $Y=3.33
+ $X2=11.28 $Y2=3.33
r215 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.48 $Y=3.33
+ $X2=11.645 $Y2=3.33
r216 71 112 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=11.81 $Y=3.33
+ $X2=12.24 $Y2=3.33
r217 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.81 $Y=3.33
+ $X2=11.645 $Y2=3.33
r218 69 105 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=3.33
+ $X2=10.32 $Y2=3.33
r219 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.485 $Y=3.33
+ $X2=10.61 $Y2=3.33
r220 68 108 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=10.735 $Y=3.33
+ $X2=11.28 $Y2=3.33
r221 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.735 $Y=3.33
+ $X2=10.61 $Y2=3.33
r222 66 91 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r223 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r224 65 95 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r225 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r226 61 64 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.705 $Y=1.985
+ $X2=12.705 $Y2=2.815
r227 59 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.705 $Y=3.245
+ $X2=12.705 $Y2=3.33
r228 59 64 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.705 $Y=3.245
+ $X2=12.705 $Y2=2.815
r229 55 58 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=11.645 $Y=2.265
+ $X2=11.645 $Y2=2.815
r230 53 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.645 $Y=3.245
+ $X2=11.645 $Y2=3.33
r231 53 58 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.645 $Y=3.245
+ $X2=11.645 $Y2=2.815
r232 49 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.61 $Y=3.245
+ $X2=10.61 $Y2=3.33
r233 49 51 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=10.61 $Y=3.245
+ $X2=10.61 $Y2=2.75
r234 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.47 $Y=1.91
+ $X2=8.47 $Y2=2.59
r235 43 129 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.47 $Y=3.245
+ $X2=8.47 $Y2=3.33
r236 43 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.47 $Y=3.245
+ $X2=8.47 $Y2=2.59
r237 42 126 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.54 $Y=3.33
+ $X2=7.372 $Y2=3.33
r238 41 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.385 $Y=3.33
+ $X2=8.47 $Y2=3.33
r239 41 42 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.385 $Y=3.33
+ $X2=7.54 $Y2=3.33
r240 37 126 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.372 $Y=3.245
+ $X2=7.372 $Y2=3.33
r241 37 39 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.372 $Y=3.245
+ $X2=7.372 $Y2=2.825
r242 33 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r243 33 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.815
r244 29 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r245 29 31 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.79
r246 25 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r247 25 27 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.465
r248 8 64 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=12.56
+ $Y=1.84 $X2=12.705 $Y2=2.815
r249 8 61 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.56
+ $Y=1.84 $X2=12.705 $Y2=1.985
r250 7 58 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=11.41
+ $Y=2.54 $X2=11.645 $Y2=2.815
r251 7 55 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=11.41
+ $Y=2.54 $X2=11.645 $Y2=2.265
r252 6 51 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=10.385
+ $Y=2.54 $X2=10.57 $Y2=2.75
r253 5 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=1.735 $X2=8.47 $Y2=2.59
r254 5 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=1.735 $X2=8.47 $Y2=1.91
r255 4 39 600 $w=1.7e-07 $l=6.26578e-07 $layer=licon1_PDIFF $count=1 $X=7.135
+ $Y=2.305 $X2=7.37 $Y2=2.825
r256 3 35 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.84 $X2=4.87 $Y2=2.815
r257 2 31 600 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.32 $X2=3.26 $Y2=2.79
r258 1 27 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.32 $X2=0.78 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%A_300_464# 1 2 3 4 5 16 20 22 25 28 29 32
+ 35 36 37 38 39 41 44 46 52
c151 38 0 1.29298e-19 $X=6.37 $Y=2.13
c152 36 0 1.57288e-19 $X=6.37 $Y=1.285
c153 32 0 6.15336e-20 $X=5.875 $Y=0.81
c154 25 0 1.19423e-19 $X=3.53 $Y=2.33
r155 50 52 17.2642 $w=2.12e-07 $l=3e-07 $layer=LI1_cond $X=3.53 $Y=2.445
+ $X2=3.83 $Y2=2.445
r156 46 48 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.435 $Y=0.68
+ $X2=2.435 $Y2=1.005
r157 43 44 10.3843 $w=6.33e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=2.662
+ $X2=2.555 $Y2=2.662
r158 40 41 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.455 $Y=1.37
+ $X2=6.455 $Y2=2.045
r159 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.37 $Y=2.13
+ $X2=6.455 $Y2=2.045
r160 38 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.37 $Y=2.13
+ $X2=6.075 $Y2=2.13
r161 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.37 $Y=1.285
+ $X2=6.455 $Y2=1.37
r162 36 37 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.37 $Y=1.285
+ $X2=5.96 $Y2=1.285
r163 35 54 3.18959 $w=2.5e-07 $l=1.67e-07 $layer=LI1_cond $X=5.95 $Y=2.39
+ $X2=5.95 $Y2=2.557
r164 34 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=6.075 $Y2=2.13
r165 34 35 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=5.95 $Y2=2.39
r166 30 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.875 $Y=1.2
+ $X2=5.96 $Y2=1.285
r167 30 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.875 $Y=1.2
+ $X2=5.875 $Y2=0.81
r168 29 52 10.0094 $w=2.12e-07 $l=1.79374e-07 $layer=LI1_cond $X=3.995 $Y=2.475
+ $X2=3.83 $Y2=2.445
r169 28 54 3.95357 $w=1.7e-07 $l=1.60857e-07 $layer=LI1_cond $X=5.825 $Y=2.475
+ $X2=5.95 $Y2=2.557
r170 28 29 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=5.825 $Y=2.475
+ $X2=3.995 $Y2=2.475
r171 25 50 2.03271 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.53 $Y=2.33
+ $X2=3.53 $Y2=2.445
r172 24 25 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.53 $Y=1.09
+ $X2=3.53 $Y2=2.33
r173 23 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=1.005
+ $X2=2.435 $Y2=1.005
r174 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=3.53 $Y2=1.09
r175 22 23 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=2.6 $Y2=1.005
r176 20 50 5.40561 $w=2.12e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=3.53 $Y2=2.445
r177 20 44 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=2.555 $Y2=2.43
r178 16 43 2.86305 $w=6.33e-07 $l=1.52e-07 $layer=LI1_cond $X=2.238 $Y=2.662
+ $X2=2.39 $Y2=2.662
r179 16 18 11.0755 $w=6.33e-07 $l=5.88e-07 $layer=LI1_cond $X=2.238 $Y=2.662
+ $X2=1.65 $Y2=2.662
r180 5 54 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.285 $X2=5.91 $Y2=2.495
r181 4 52 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.68
+ $Y=2.32 $X2=3.83 $Y2=2.465
r182 3 43 200 $w=1.7e-07 $l=9.59766e-07 $layer=licon1_PDIFF $count=3 $X=1.5
+ $Y=2.32 $X2=2.39 $Y2=2.465
r183 3 18 200 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=3 $X=1.5
+ $Y=2.32 $X2=1.65 $Y2=2.465
r184 2 32 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=5.73
+ $Y=0.59 $X2=5.875 $Y2=0.81
r185 1 46 182 $w=1.7e-07 $l=6.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.405 $X2=2.435 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%Q 1 2 7 8 9 10 11 12 13 29
r15 22 29 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=13.16 $Y=0.965
+ $X2=13.16 $Y2=0.925
r16 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=13.197 $Y=2.405
+ $X2=13.197 $Y2=2.775
r17 11 12 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=13.197 $Y=1.985
+ $X2=13.197 $Y2=2.405
r18 10 11 14.462 $w=2.53e-07 $l=3.2e-07 $layer=LI1_cond $X=13.197 $Y=1.665
+ $X2=13.197 $Y2=1.985
r19 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=13.197 $Y=1.295
+ $X2=13.197 $Y2=1.665
r20 9 45 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=13.197 $Y=1.295
+ $X2=13.197 $Y2=1.13
r21 8 45 5.6192 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=13.16 $Y=0.987
+ $X2=13.16 $Y2=1.13
r22 8 22 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=13.16 $Y=0.987
+ $X2=13.16 $Y2=0.965
r23 8 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=13.16 $Y=0.902
+ $X2=13.16 $Y2=0.925
r24 7 8 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=13.16 $Y=0.515
+ $X2=13.16 $Y2=0.902
r25 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=1.84 $X2=13.155 $Y2=2.815
r26 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=1.84 $X2=13.155 $Y2=1.985
r27 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.02
+ $Y=0.37 $X2=13.16 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 47 48
+ 50 51 52 54 69 73 81 86 93 94 97 101 107 110 113
c126 94 0 7.12888e-20 $X=13.2 $Y=0
c127 32 0 6.15093e-20 $X=4.88 $Y=0.55
r128 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r129 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r130 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r131 101 104 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.595 $Y2=0.325
r132 101 102 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r133 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r134 94 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r135 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r136 91 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.815 $Y=0
+ $X2=12.69 $Y2=0
r137 91 93 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.815 $Y=0
+ $X2=13.2 $Y2=0
r138 90 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r139 90 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r140 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r141 87 110 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=11.737 $Y2=0
r142 87 89 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=12.24 $Y2=0
r143 86 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.565 $Y=0
+ $X2=12.69 $Y2=0
r144 86 89 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.565 $Y=0
+ $X2=12.24 $Y2=0
r145 85 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r146 85 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r147 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r148 82 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.525 $Y=0
+ $X2=10.36 $Y2=0
r149 82 84 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=10.525 $Y=0
+ $X2=11.28 $Y2=0
r150 81 110 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=11.57 $Y=0
+ $X2=11.737 $Y2=0
r151 81 84 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=11.57 $Y=0
+ $X2=11.28 $Y2=0
r152 80 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r153 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r154 77 80 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r155 77 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r156 76 79 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r157 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r158 74 101 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.595 $Y2=0
r159 74 76 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.92
+ $Y2=0
r160 73 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=10.36 $Y2=0
r161 73 79 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=9.84 $Y2=0
r162 71 72 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r163 69 101 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=7.595 $Y2=0
r164 69 71 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=7.43 $Y=0 $X2=5.04
+ $Y2=0
r165 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r166 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r167 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r168 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r169 62 65 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r170 62 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r171 61 64 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r172 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r173 59 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r174 59 61 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r175 57 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r176 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r177 54 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r178 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r179 52 102 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=7.44 $Y2=0
r180 52 72 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=5.04 $Y2=0
r181 50 67 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=4.56 $Y2=0
r182 50 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.84
+ $Y2=0
r183 49 71 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.965 $Y=0 $X2=5.04
+ $Y2=0
r184 49 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.965 $Y=0 $X2=4.84
+ $Y2=0
r185 47 64 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.6
+ $Y2=0
r186 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.87
+ $Y2=0
r187 46 67 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=4.56 $Y2=0
r188 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.87
+ $Y2=0
r189 42 113 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.69 $Y=0.085
+ $X2=12.69 $Y2=0
r190 42 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.69 $Y=0.085
+ $X2=12.69 $Y2=0.515
r191 38 110 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=11.737 $Y=0.085
+ $X2=11.737 $Y2=0
r192 38 40 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=11.737 $Y=0.085
+ $X2=11.737 $Y2=0.5
r193 34 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0
r194 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0.58
r195 30 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0
r196 30 32 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0.55
r197 26 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0.085
+ $X2=3.87 $Y2=0
r198 26 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.87 $Y=0.085
+ $X2=3.87 $Y2=0.565
r199 22 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r200 22 24 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.65
r201 7 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.585
+ $Y=0.37 $X2=12.73 $Y2=0.515
r202 6 40 182 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=1 $X=11.59
+ $Y=0.37 $X2=11.735 $Y2=0.5
r203 5 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.22
+ $Y=0.37 $X2=10.36 $Y2=0.58
r204 4 104 182 $w=1.7e-07 $l=3.58504e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.59 $X2=7.595 $Y2=0.325
r205 3 32 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.74 $Y=0.37
+ $X2=4.88 $Y2=0.55
r206 2 28 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.405 $X2=3.87 $Y2=0.565
r207 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.44 $X2=0.71 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_1%noxref_24 1 2 7 9
c25 7 0 8.6114e-20 $X=3.09 $Y=0.34
r26 9 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=0.34 $X2=1.27
+ $Y2=0.55
r27 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34 $X2=1.27
+ $Y2=0.34
r28 7 17 4.87721 $w=5.13e-07 $l=2.1e-07 $layer=LI1_cond $X=3.347 $Y=0.34
+ $X2=3.347 $Y2=0.55
r29 7 8 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=3.09 $Y=0.34
+ $X2=1.435 $Y2=0.34
r30 2 17 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.405 $X2=3.345 $Y2=0.55
r31 1 12 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.55
.ends

