* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1827_144# a_1074_88# a_1429_308# VPB pshort w=1e+06u l=150000u
+  ad=3.128e+11p pd=2.73e+06u as=7.85e+11p ps=3.57e+06u
M1001 VGND a_2087_410# a_2073_74# VNB nlowvt w=420000u l=150000u
+  ad=1.79055e+12p pd=1.44e+07u as=1.05e+11p ps=1.34e+06u
M1002 a_284_464# D a_206_464# VPB pshort w=640000u l=150000u
+  ad=8.151e+11p pd=6.15e+06u as=1.536e+11p ps=1.76e+06u
M1003 a_538_81# SCE a_284_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.549e+11p ps=3.37e+06u
M1004 a_2265_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1005 a_2087_410# a_1827_144# a_2265_74# VNB nlowvt w=420000u l=150000u
+  ad=2.1e+11p pd=1.84e+06u as=0p ps=0u
M1006 VPWR SCD a_471_464# VPB pshort w=640000u l=150000u
+  ad=2.58055e+12p pd=2.111e+07u as=1.536e+11p ps=1.76e+06u
M1007 VPWR a_1429_308# a_1384_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 VPWR a_1827_144# a_2492_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 a_854_74# CLK_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 Q a_2492_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1011 a_1272_131# RESET_B VPWR VPB pshort w=420000u l=150000u
+  ad=2.499e+11p pd=2.87e+06u as=0p ps=0u
M1012 a_284_464# RESET_B VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_324_81# a_27_88# a_239_81# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.373e+11p ps=2.81e+06u
M1014 a_284_464# D a_324_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1074_88# a_854_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 VPWR SCE a_27_88# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1017 a_206_464# SCE VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND RESET_B a_1489_131# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 Q a_2492_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1020 a_1272_131# a_854_74# a_284_464# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_2087_410# a_2042_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1022 VGND RESET_B a_239_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1411_131# a_854_74# a_1272_131# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.289e+11p ps=1.93e+06u
M1024 a_1384_508# a_1074_88# a_1272_131# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1429_308# a_1272_131# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1074_88# a_854_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1027 a_1272_131# a_1074_88# a_284_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_2073_74# a_1074_88# a_1827_144# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=6.2565e+11p ps=4.26e+06u
M1029 VGND a_1827_144# a_2492_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1030 a_2087_410# RESET_B VPWR VPB pshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1031 a_2042_508# a_854_74# a_1827_144# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_1827_144# a_2087_410# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_239_81# SCD a_538_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1489_131# a_1429_308# a_1411_131# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1429_308# a_1272_131# VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=2.4e+06u as=0p ps=0u
M1036 a_471_464# a_27_88# a_284_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND SCE a_27_88# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1038 a_854_74# CLK_N VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1039 a_1827_144# a_854_74# a_1429_308# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
