* File: sky130_fd_sc_hs__nand3_2.pex.spice
* Created: Tue Sep  1 20:09:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND3_2%C 1 3 4 6 7 9 10 12 13 19 20
c51 20 0 1.06079e-19 $X=0.91 $Y=1.492
c52 19 0 6.03852e-20 $X=0.57 $Y=1.385
c53 10 0 1.8621e-19 $X=0.955 $Y=1.765
r54 20 21 4.98621 $w=4.35e-07 $l=4.5e-08 $layer=POLY_cond $X=0.91 $Y=1.492
+ $X2=0.955 $Y2=1.492
r55 18 20 37.6736 $w=4.35e-07 $l=3.4e-07 $layer=POLY_cond $X=0.57 $Y=1.492
+ $X2=0.91 $Y2=1.492
r56 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.57
+ $Y=1.385 $X2=0.57 $Y2=1.385
r57 16 18 7.2023 $w=4.35e-07 $l=6.5e-08 $layer=POLY_cond $X=0.505 $Y=1.492
+ $X2=0.57 $Y2=1.492
r58 15 16 2.77011 $w=4.35e-07 $l=2.5e-08 $layer=POLY_cond $X=0.48 $Y=1.492
+ $X2=0.505 $Y2=1.492
r59 13 19 10.2785 $w=3.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.57 $Y2=1.365
r60 10 21 27.9254 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.492
r61 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r62 7 20 27.9254 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.91 $Y=1.22
+ $X2=0.91 $Y2=1.492
r63 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.91 $Y=1.22 $X2=0.91
+ $Y2=0.74
r64 4 16 27.9254 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.492
r65 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r66 1 15 27.9254 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.48 $Y=1.22
+ $X2=0.48 $Y2=1.492
r67 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.48 $Y=1.22 $X2=0.48
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_2%B 3 5 7 8 10 13 15 16 18 23 26 33 38
c92 26 0 9.2975e-20 $X=1.595 $Y=1.58
c93 16 0 1.8621e-19 $X=1.795 $Y=2.035
c94 5 0 1.34415e-19 $X=1.455 $Y=1.765
c95 3 0 6.03852e-20 $X=1.34 $Y=0.74
r96 33 38 0.721711 $w=4.34e-07 $l=8.7178e-08 $layer=LI1_cond $X=1.61 $Y=1.68
+ $X2=1.53 $Y2=1.665
r97 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.515 $X2=1.43 $Y2=1.515
r98 26 38 0.983871 $w=4.34e-07 $l=3.5e-08 $layer=LI1_cond $X=1.53 $Y=1.63
+ $X2=1.53 $Y2=1.665
r99 26 31 3.23272 $w=4.34e-07 $l=1.15e-07 $layer=LI1_cond $X=1.53 $Y=1.63
+ $X2=1.53 $Y2=1.515
r100 26 33 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.61 $Y=1.715
+ $X2=1.61 $Y2=1.68
r101 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.9
+ $Y=1.485 $X2=2.9 $Y2=1.485
r102 20 23 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.74 $Y=1.485
+ $X2=2.9 $Y2=1.485
r103 19 26 7.31957 $w=3.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.61 $Y=1.95
+ $X2=1.61 $Y2=1.715
r104 17 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=1.65
+ $X2=2.74 $Y2=1.485
r105 17 18 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.74 $Y=1.65 $X2=2.74
+ $Y2=1.95
r106 16 19 8.10976 $w=1.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.795 $Y=2.035
+ $X2=1.61 $Y2=1.95
r107 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.655 $Y=2.035
+ $X2=2.74 $Y2=1.95
r108 15 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.655 $Y=2.035
+ $X2=1.795 $Y2=2.035
r109 11 24 38.6072 $w=2.91e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.88 $Y=1.32
+ $X2=2.9 $Y2=1.485
r110 11 13 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.88 $Y=1.32
+ $X2=2.88 $Y2=0.795
r111 8 24 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.9 $Y2=1.485
r112 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r113 5 30 52.2586 $w=2.99e-07 $l=2.62202e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.43 $Y2=1.515
r114 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r115 1 30 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.34 $Y=1.35
+ $X2=1.43 $Y2=1.515
r116 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.34 $Y=1.35 $X2=1.34
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_2%A 3 5 7 10 12 14 15 21 22
c57 10 0 5.74086e-20 $X=2.325 $Y=0.795
r58 22 23 10.2827 $w=3.75e-07 $l=8e-08 $layer=POLY_cond $X=2.325 $Y=1.557
+ $X2=2.405 $Y2=1.557
r59 20 22 25.064 $w=3.75e-07 $l=1.95e-07 $layer=POLY_cond $X=2.13 $Y=1.557
+ $X2=2.325 $Y2=1.557
r60 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r61 18 20 28.2773 $w=3.75e-07 $l=2.2e-07 $layer=POLY_cond $X=1.91 $Y=1.557
+ $X2=2.13 $Y2=1.557
r62 17 18 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=1.895 $Y=1.557
+ $X2=1.91 $Y2=1.557
r63 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.515
r64 12 23 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.557
r65 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r66 8 22 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.325 $Y=1.35
+ $X2=2.325 $Y2=1.557
r67 8 10 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.325 $Y=1.35
+ $X2=2.325 $Y2=0.795
r68 5 18 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=1.557
r69 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=2.4
r70 1 17 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.895 $Y=1.35
+ $X2=1.895 $Y2=1.557
r71 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.895 $Y=1.35
+ $X2=1.895 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_2%VPWR 1 2 3 4 13 15 21 25 27 29 33 35 40 45
+ 54 57 61
r57 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 49 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 49 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 46 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.18 $Y2=3.33
r65 46 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 45 60 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.177 $Y2=3.33
r67 45 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 41 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.19 $Y2=3.33
r69 41 43 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 40 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.18 $Y2=3.33
r71 40 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 36 51 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r76 36 38 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 35 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.19 $Y2=3.33
r78 35 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 33 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r80 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r81 33 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r82 29 32 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.12 $Y=1.985
+ $X2=3.12 $Y2=2.815
r83 27 60 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.177 $Y2=3.33
r84 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=2.815
r85 23 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=3.33
r86 23 25 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=2.795
r87 19 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=3.33
r88 19 21 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.795
r89 15 18 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r90 13 51 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r91 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r92 4 32 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.815
r93 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=1.985
r94 3 25 600 $w=1.7e-07 $l=1.04797e-06 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.18 $Y2=2.795
r95 2 21 600 $w=1.7e-07 $l=1.05025e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.795
r96 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r97 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_2%Y 1 2 3 4 15 19 20 21 23 25 27 30 31 35 41
+ 42
c87 30 0 1.34415e-19 $X=0.73 $Y=1.985
c88 19 0 5.74086e-20 $X=1.945 $Y=1.175
r89 41 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.375
+ $X2=1.68 $Y2=2.46
r90 41 42 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=2.475 $X2=1.68
+ $Y2=2.775
r91 41 46 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.68 $Y=2.475
+ $X2=1.68 $Y2=2.46
r92 35 37 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.11 $Y=1.02
+ $X2=2.11 $Y2=1.175
r93 32 33 3.61166 $w=5.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=2.375
+ $X2=0.83 $Y2=2.46
r94 30 32 8.80133 $w=5.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.83 $Y=1.985
+ $X2=0.83 $Y2=2.375
r95 30 31 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.83 $Y=1.985
+ $X2=0.83 $Y2=1.82
r96 25 40 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.46 $X2=2.66
+ $Y2=2.375
r97 25 27 15.1525 $w=2.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.66 $Y=2.46
+ $X2=2.66 $Y2=2.815
r98 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.375
+ $X2=1.68 $Y2=2.375
r99 23 40 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=2.375
+ $X2=2.66 $Y2=2.375
r100 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.525 $Y=2.375
+ $X2=1.845 $Y2=2.375
r101 22 32 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.095 $Y=2.375
+ $X2=0.83 $Y2=2.375
r102 21 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.375
+ $X2=1.68 $Y2=2.375
r103 21 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.515 $Y=2.375
+ $X2=1.095 $Y2=2.375
r104 19 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=1.175
+ $X2=2.11 $Y2=1.175
r105 19 20 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.945 $Y=1.175
+ $X2=1.095 $Y2=1.175
r106 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.01 $Y=1.26
+ $X2=1.095 $Y2=1.175
r107 17 31 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.01 $Y=1.26
+ $X2=1.01 $Y2=1.82
r108 15 33 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.73 $Y=2.815
+ $X2=0.73 $Y2=2.46
r109 4 40 600 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.375
r110 4 27 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.815
r111 3 41 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.41
r112 2 30 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r113 2 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r114 1 35 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.425 $X2=2.11 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_2%A_27_74# 1 2 3 12 14 16 20 27 30
c59 27 0 1.31036e-20 $X=1.205 $Y=0.68
r60 27 28 7.32946 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=1.205 $Y=0.68
+ $X2=1.205 $Y2=0.835
r61 26 27 8.74806 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=1.205 $Y=0.495
+ $X2=1.205 $Y2=0.68
r62 20 23 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=0.265 $Y=0.835
+ $X2=0.265 $Y2=0.895
r63 20 21 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=0.835
+ $X2=0.265 $Y2=0.75
r64 17 27 3.17874 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=0.68
+ $X2=1.205 $Y2=0.68
r65 16 30 4.5891 $w=1.7e-07 $l=2.07123e-07 $layer=LI1_cond $X=2.93 $Y=0.68
+ $X2=3.095 $Y2=0.585
r66 16 17 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=2.93 $Y=0.68
+ $X2=1.37 $Y2=0.68
r67 15 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.43 $Y=0.835
+ $X2=0.265 $Y2=0.835
r68 14 28 3.17874 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=0.835
+ $X2=1.205 $Y2=0.835
r69 14 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.04 $Y=0.835
+ $X2=0.43 $Y2=0.835
r70 12 21 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=0.225 $Y=0.515
+ $X2=0.225 $Y2=0.75
r71 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.955
+ $Y=0.425 $X2=3.095 $Y2=0.57
r72 2 26 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.37 $X2=1.125 $Y2=0.495
r73 1 23 182 $w=1.7e-07 $l=5.86409e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.265 $Y2=0.895
r74 1 12 182 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_2%VGND 1 6 8 10 20 21 24
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 17 20 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r44 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=0.695
+ $Y2=0
r46 15 17 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=1.2
+ $Y2=0
r47 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r48 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r49 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.695
+ $Y2=0
r50 10 12 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.24
+ $Y2=0
r51 8 21 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r52 8 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r53 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r54 4 6 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.495
r55 1 6 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.37 $X2=0.695 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_2%A_283_74# 1 2 11
r16 8 11 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=1.62 $Y=0.34 $X2=2.6
+ $Y2=0.34
r17 2 11 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.425 $X2=2.6 $Y2=0.34
r18 1 8 182 $w=1.7e-07 $l=2.19488e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.37 $X2=1.62 $Y2=0.34
.ends

