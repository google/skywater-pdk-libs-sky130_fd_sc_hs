* File: sky130_fd_sc_hs__a22oi_4.spice
* Created: Thu Aug 27 20:27:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a22oi_4.pex.spice"
.subckt sky130_fd_sc_hs__a22oi_4  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_B2_M1008_g N_A_48_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1008_d N_B2_M1013_g N_A_48_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_B2_M1016_g N_A_48_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1016_d N_B2_M1025_g N_A_48_74#_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1004 N_A_48_74#_M1025_s N_B1_M1004_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1005 N_A_48_74#_M1005_d N_B1_M1005_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1021 N_A_48_74#_M1005_d N_B1_M1021_g N_Y_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_A_48_74#_M1022_d N_B1_M1022_g N_Y_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_840_74#_M1012_d N_A1_M1012_g N_Y_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1018 N_A_840_74#_M1018_d N_A1_M1018_g N_Y_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1024 N_A_840_74#_M1018_d N_A1_M1024_g N_Y_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1029 N_A_840_74#_M1029_d N_A1_M1029_g N_Y_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A2_M1014_g N_A_840_74#_M1029_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1014_d N_A2_M1015_g N_A_840_74#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A2_M1017_g N_A_840_74#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1017_d N_A2_M1028_g N_A_840_74#_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_Y_M1019_d N_B2_M1019_g N_A_45_368#_M1019_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007.2 A=0.168 P=2.54 MULT=1
MM1023 N_Y_M1019_d N_B2_M1023_g N_A_45_368#_M1023_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75006.7 A=0.168 P=2.54 MULT=1
MM1026 N_Y_M1026_d N_B2_M1026_g N_A_45_368#_M1023_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75006.3 A=0.168 P=2.54 MULT=1
MM1030 N_Y_M1026_d N_B2_M1030_g N_A_45_368#_M1030_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75005.8 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_45_368#_M1030_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75005.4 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1001_d N_B1_M1002_g N_A_45_368#_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_A_45_368#_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75004.5 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1006_d N_B1_M1007_g N_A_45_368#_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75004 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_45_368#_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.8 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1010_d N_A1_M1011_g N_A_45_368#_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.2 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1020 N_VPWR_M1020_d N_A1_M1020_g N_A_45_368#_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2968 AS=0.168 PD=1.65 PS=1.42 NRD=21.9852 NRS=1.7533 M=1 R=7.46667
+ SA=75004.7 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1027 N_VPWR_M1020_d N_A1_M1027_g N_A_45_368#_M1027_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2968 AS=0.168 PD=1.65 PS=1.42 NRD=21.9852 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75002 A=0.168 P=2.54 MULT=1
MM1000 N_A_45_368#_M1027_s N_A2_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.8 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1003 N_A_45_368#_M1003_d N_A2_M1003_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.3 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1009 N_A_45_368#_M1003_d N_A2_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.7 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1031 N_A_45_368#_M1031_d N_A2_M1031_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_hs__a22oi_4.pxi.spice"
*
.ends
*
*
