* NGSPICE file created from sky130_fd_sc_hs__a221oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_118_368# C1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=6.44e+11p pd=5.63e+06u as=3.08e+11p ps=2.79e+06u
M1001 Y B1 a_351_74# VNB nlowvt w=740000u l=150000u
+  ad=8.695e+11p pd=5.31e+06u as=1.554e+11p ps=1.9e+06u
M1002 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=0p ps=0u
M1003 a_567_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1004 VGND A2 a_567_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_118_368# B2 a_263_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=9.856e+11p ps=8.48e+06u
M1006 VPWR A1 a_263_368# VPB pshort w=1.12e+06u l=150000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1007 a_351_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_263_368# B1 a_118_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_263_368# A2 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

