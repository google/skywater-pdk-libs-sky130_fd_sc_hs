* File: sky130_fd_sc_hs__o311a_2.spice
* Created: Thu Aug 27 21:01:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o311a_2.pex.spice"
.subckt sky130_fd_sc_hs__o311a_2  VNB VPB C1 B1 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1001 A_135_74# N_C1_M1001_g N_A_32_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0999 AS=0.2701 PD=1.01 PS=2.21 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1012 N_A_219_74#_M1012_d N_B1_M1012_g A_135_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.0999 PD=1.13 PS=1.01 NRD=17.832 NRS=12.972 M=1 R=4.93333
+ SA=75000.7 SB=75003 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A3_M1004_g N_A_219_74#_M1012_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2487 AS=0.1443 PD=1.49 PS=1.13 NRD=45.576 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1000 N_A_219_74#_M1000_d N_A2_M1000_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2487 PD=1.02 PS=1.49 NRD=0 NRS=45.576 M=1 R=4.93333 SA=75002
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A1_M1008_g N_A_219_74#_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.16465 AS=0.1036 PD=1.185 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1006 N_X_M1006_d N_A_32_74#_M1006_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.16465 PD=1.02 PS=1.185 NRD=0 NRS=15.396 M=1 R=4.93333 SA=75003
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1006_d N_A_32_74#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2775 PD=1.02 PS=2.23 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75003.4
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_C1_M1010_g N_A_32_74#_M1010_s VPB PSHORT L=0.15 W=1
+ AD=0.21 AS=0.295 PD=1.42 PS=2.59 NRD=21.67 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1013 N_A_32_74#_M1013_d N_B1_M1013_g N_VPWR_M1010_d VPB PSHORT L=0.15 W=1
+ AD=0.20066 AS=0.21 PD=1.42453 PS=1.42 NRD=20.0152 NRS=5.8903 M=1 R=6.66667
+ SA=75000.8 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1005 A_360_368# N_A3_M1005_g N_A_32_74#_M1013_d VPB PSHORT L=0.15 W=1.12
+ AD=0.1512 AS=0.22474 PD=1.39 PS=1.59547 NRD=14.0658 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1007 A_444_368# N_A2_M1007_g A_360_368# VPB PSHORT L=0.15 W=1.12 AD=0.2184
+ AS=0.1512 PD=1.51 PS=1.39 NRD=24.6053 NRS=14.0658 M=1 R=7.46667 SA=75001.6
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g A_444_368# VPB PSHORT L=0.15 W=1.12 AD=0.2436
+ AS=0.2184 PD=1.555 PS=1.51 NRD=1.7533 NRS=24.6053 M=1 R=7.46667 SA=75002.2
+ SB=75001.3 A=0.168 P=2.54 MULT=1
MM1002 N_X_M1002_d N_A_32_74#_M1002_g N_VPWR_M1011_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2436 PD=1.42 PS=1.555 NRD=1.7533 NRS=25.4918 M=1 R=7.46667
+ SA=75002.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1003 N_X_M1002_d N_A_32_74#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.2 SB=75000.3 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__o311a_2.pxi.spice"
*
.ends
*
*
