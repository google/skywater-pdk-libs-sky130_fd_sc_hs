* File: sky130_fd_sc_hs__a311oi_1.pxi.spice
* Created: Tue Sep  1 19:52:32 2020
* 
x_PM_SKY130_FD_SC_HS__A311OI_1%A3 N_A3_c_60_n N_A3_M1000_g N_A3_M1004_g
+ N_A3_c_57_n N_A3_c_58_n A3 A3 PM_SKY130_FD_SC_HS__A311OI_1%A3
x_PM_SKY130_FD_SC_HS__A311OI_1%A2 N_A2_M1002_g N_A2_c_85_n N_A2_M1001_g A2
+ N_A2_c_86_n PM_SKY130_FD_SC_HS__A311OI_1%A2
x_PM_SKY130_FD_SC_HS__A311OI_1%A1 N_A1_M1006_g N_A1_c_117_n N_A1_M1007_g A1
+ N_A1_c_118_n PM_SKY130_FD_SC_HS__A311OI_1%A1
x_PM_SKY130_FD_SC_HS__A311OI_1%B1 N_B1_M1009_g N_B1_c_146_n N_B1_M1008_g B1 B1
+ PM_SKY130_FD_SC_HS__A311OI_1%B1
x_PM_SKY130_FD_SC_HS__A311OI_1%C1 N_C1_M1003_g N_C1_c_179_n N_C1_M1005_g
+ N_C1_c_176_n C1 N_C1_c_177_n N_C1_c_178_n PM_SKY130_FD_SC_HS__A311OI_1%C1
x_PM_SKY130_FD_SC_HS__A311OI_1%VPWR N_VPWR_M1000_s N_VPWR_M1001_d N_VPWR_c_206_n
+ N_VPWR_c_207_n N_VPWR_c_208_n N_VPWR_c_209_n N_VPWR_c_210_n N_VPWR_c_211_n
+ VPWR N_VPWR_c_212_n N_VPWR_c_205_n PM_SKY130_FD_SC_HS__A311OI_1%VPWR
x_PM_SKY130_FD_SC_HS__A311OI_1%A_156_368# N_A_156_368#_M1000_d
+ N_A_156_368#_M1007_d N_A_156_368#_c_243_n N_A_156_368#_c_240_n
+ N_A_156_368#_c_241_n PM_SKY130_FD_SC_HS__A311OI_1%A_156_368#
x_PM_SKY130_FD_SC_HS__A311OI_1%Y N_Y_M1006_d N_Y_M1003_d N_Y_M1005_d N_Y_c_268_n
+ N_Y_c_280_n N_Y_c_286_n N_Y_c_281_n N_Y_c_269_n N_Y_c_270_n N_Y_c_274_n
+ N_Y_c_275_n Y Y N_Y_c_271_n N_Y_c_272_n PM_SKY130_FD_SC_HS__A311OI_1%Y
x_PM_SKY130_FD_SC_HS__A311OI_1%VGND N_VGND_M1004_s N_VGND_M1009_d N_VGND_c_337_n
+ N_VGND_c_338_n N_VGND_c_339_n N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n
+ VGND N_VGND_c_343_n N_VGND_c_344_n PM_SKY130_FD_SC_HS__A311OI_1%VGND
cc_1 VNB N_A3_c_57_n 0.0696532f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_2 VNB N_A3_c_58_n 0.0197654f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.22
cc_3 VNB A3 0.0295507f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A2_M1002_g 0.0244269f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_5 VNB N_A2_c_85_n 0.0262555f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_6 VNB N_A2_c_86_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A1_M1006_g 0.0268314f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_8 VNB N_A1_c_117_n 0.0262348f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_9 VNB N_A1_c_118_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_M1009_g 0.0261863f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_11 VNB N_B1_c_146_n 0.0216541f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_12 VNB B1 0.00423229f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.22
cc_13 VNB N_C1_M1003_g 0.0345407f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_14 VNB N_C1_c_176_n 0.00982321f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.22
cc_15 VNB N_C1_c_177_n 0.0439496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_c_178_n 0.00813406f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.385
cc_17 VNB N_VPWR_c_205_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_268_n 0.00348446f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_Y_c_269_n 0.0134556f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.385
cc_20 VNB N_Y_c_270_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_271_n 0.00580575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_272_n 0.0242391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_337_n 0.0285265f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.22
cc_24 VNB N_VGND_c_338_n 0.00685406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_339_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.385
cc_26 VNB N_VGND_c_340_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_341_n 0.0411805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_342_n 0.0069273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_343_n 0.0244021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_344_n 0.225214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_A3_c_60_n 0.0177645f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_32 VPB N_A3_c_57_n 0.00686864f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.385
cc_33 VPB A3 0.0162112f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_34 VPB N_A2_c_85_n 0.0279855f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_35 VPB N_A2_c_86_n 0.00299909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A1_c_117_n 0.0284701f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_37 VPB N_A1_c_118_n 0.00244477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_B1_c_146_n 0.0265378f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_39 VPB B1 0.00488575f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.22
cc_40 VPB N_C1_c_179_n 0.021323f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_41 VPB N_C1_c_176_n 0.00609676f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.22
cc_42 VPB N_C1_c_177_n 0.0145157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_C1_c_178_n 0.0117196f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_44 VPB N_VPWR_c_206_n 0.0380055f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.22
cc_45 VPB N_VPWR_c_207_n 0.0106054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_208_n 0.0121672f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_47 VPB N_VPWR_c_209_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_210_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_211_n 0.00786036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_212_n 0.0506387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_205_n 0.0850486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_156_368#_c_240_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_53 VPB N_A_156_368#_c_241_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_54 VPB N_Y_c_268_n 0.00133931f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_55 VPB N_Y_c_274_n 0.00743317f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_56 VPB N_Y_c_275_n 0.0360166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 N_A3_c_58_n N_A2_M1002_g 0.0431169f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A3_c_60_n N_A2_c_85_n 0.0242467f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_59 N_A3_c_57_n N_A2_c_85_n 0.0471303f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_60 N_A3_c_57_n N_A2_c_86_n 6.49042e-19 $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_61 N_A3_c_60_n N_VPWR_c_206_n 0.0071424f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_62 A3 N_VPWR_c_206_n 0.00741364f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A3_c_60_n N_VPWR_c_210_n 0.00445602f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A3_c_60_n N_VPWR_c_205_n 0.00861667f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A3_c_60_n N_A_156_368#_c_240_n 0.00815828f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_66 N_A3_c_60_n N_Y_c_268_n 0.00923194f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_67 N_A3_c_57_n N_Y_c_268_n 0.014292f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_68 N_A3_c_58_n N_Y_c_268_n 7.61601e-19 $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_69 A3 N_Y_c_268_n 0.0442649f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A3_c_58_n N_Y_c_280_n 0.0174993f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_71 N_A3_c_60_n N_Y_c_281_n 0.0166918f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A3_c_58_n N_Y_c_272_n 0.00235309f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_73 N_A3_c_57_n N_VGND_c_337_n 0.00535484f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_74 N_A3_c_58_n N_VGND_c_337_n 0.0158743f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_75 A3 N_VGND_c_337_n 0.0085354f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A3_c_58_n N_VGND_c_341_n 0.00383152f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_77 N_A3_c_58_n N_VGND_c_344_n 0.0075694f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_78 N_A2_M1002_g N_A1_M1006_g 0.0343434f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_79 N_A2_c_85_n N_A1_c_117_n 0.0507408f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A2_c_86_n N_A1_c_117_n 0.00144235f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A2_c_85_n N_A1_c_118_n 0.0014822f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A2_c_86_n N_A1_c_118_n 0.0280928f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_83 N_A2_c_85_n N_VPWR_c_207_n 0.00591952f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A2_c_85_n N_VPWR_c_210_n 0.00445602f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A2_c_85_n N_VPWR_c_205_n 0.00858468f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A2_c_85_n N_A_156_368#_c_243_n 0.0125526f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A2_c_85_n N_A_156_368#_c_240_n 0.00783743f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A2_c_85_n N_A_156_368#_c_241_n 7.96421e-19 $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A2_M1002_g N_Y_c_268_n 0.0051053f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A2_c_85_n N_Y_c_268_n 0.00173556f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A2_c_86_n N_Y_c_268_n 0.0327278f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_92 N_A2_c_85_n N_Y_c_286_n 0.0120818f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A2_c_86_n N_Y_c_286_n 0.0210863f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A2_M1002_g N_Y_c_271_n 0.00731318f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A2_c_86_n N_Y_c_271_n 0.0268379f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A2_M1002_g N_Y_c_272_n 0.0279819f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A2_c_85_n N_Y_c_272_n 0.00140815f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A2_M1002_g N_VGND_c_337_n 0.00186934f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A2_M1002_g N_VGND_c_341_n 0.00382217f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A2_M1002_g N_VGND_c_344_n 0.00652989f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A1_M1006_g N_B1_M1009_g 0.0215861f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A1_c_117_n N_B1_c_146_n 0.0507499f $X=1.785 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A1_c_118_n N_B1_c_146_n 5.07076e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A1_c_117_n B1 0.00261368f $X=1.785 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A1_c_118_n B1 0.036282f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A1_c_117_n N_VPWR_c_207_n 0.00591952f $X=1.785 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A1_c_117_n N_VPWR_c_212_n 0.00445602f $X=1.785 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A1_c_117_n N_VPWR_c_205_n 0.00858468f $X=1.785 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A1_c_117_n N_A_156_368#_c_243_n 0.0125526f $X=1.785 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A1_c_117_n N_A_156_368#_c_240_n 7.96421e-19 $X=1.785 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A1_c_117_n N_A_156_368#_c_241_n 0.00783743f $X=1.785 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_A1_c_117_n N_Y_c_286_n 0.0121564f $X=1.785 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A1_c_118_n N_Y_c_286_n 0.0226548f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A1_M1006_g N_Y_c_272_n 0.0297967f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A1_c_117_n N_Y_c_272_n 0.0014007f $X=1.785 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A1_c_118_n N_Y_c_272_n 0.0275097f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_117 N_A1_M1006_g N_VGND_c_338_n 6.64319e-19 $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A1_M1006_g N_VGND_c_341_n 0.00291649f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A1_M1006_g N_VGND_c_344_n 0.00361179f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_120 N_B1_M1009_g N_C1_M1003_g 0.0254529f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_121 N_B1_c_146_n N_C1_c_179_n 0.0486247f $X=2.235 $Y=1.765 $X2=0 $Y2=0
cc_122 B1 N_C1_c_179_n 0.00202917f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_123 N_B1_c_146_n N_C1_c_176_n 0.0250068f $X=2.235 $Y=1.765 $X2=0 $Y2=0
cc_124 B1 N_C1_c_176_n 0.0165148f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_125 B1 N_C1_c_178_n 0.0346459f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_126 N_B1_c_146_n N_VPWR_c_212_n 0.00445602f $X=2.235 $Y=1.765 $X2=0 $Y2=0
cc_127 N_B1_c_146_n N_VPWR_c_205_n 0.00858782f $X=2.235 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B1_c_146_n N_A_156_368#_c_241_n 0.013263f $X=2.235 $Y=1.765 $X2=0 $Y2=0
cc_129 N_B1_c_146_n N_Y_c_286_n 0.0155772f $X=2.235 $Y=1.765 $X2=0 $Y2=0
cc_130 B1 N_Y_c_286_n 0.0485699f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_131 N_B1_M1009_g N_Y_c_269_n 0.0153799f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_132 N_B1_c_146_n N_Y_c_269_n 0.00434748f $X=2.235 $Y=1.765 $X2=0 $Y2=0
cc_133 B1 N_Y_c_269_n 0.0544915f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_134 N_B1_M1009_g N_Y_c_270_n 8.78222e-19 $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_135 N_B1_c_146_n N_Y_c_275_n 0.00286856f $X=2.235 $Y=1.765 $X2=0 $Y2=0
cc_136 N_B1_M1009_g N_Y_c_272_n 0.00384236f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_137 N_B1_M1009_g N_VGND_c_338_n 0.0113145f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B1_M1009_g N_VGND_c_341_n 0.00383152f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_139 N_B1_M1009_g N_VGND_c_344_n 0.00758569f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_140 N_C1_c_179_n N_VPWR_c_212_n 0.00445602f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_141 N_C1_c_179_n N_VPWR_c_205_n 0.00862572f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_142 N_C1_c_179_n N_A_156_368#_c_241_n 0.00207206f $X=2.715 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_C1_c_179_n N_Y_c_286_n 0.0126989f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_144 N_C1_M1003_g N_Y_c_269_n 0.0145657f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_145 N_C1_c_176_n N_Y_c_269_n 0.00676585f $X=2.715 $Y=1.557 $X2=0 $Y2=0
cc_146 N_C1_c_177_n N_Y_c_269_n 0.00121887f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_147 N_C1_c_178_n N_Y_c_269_n 0.0132907f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_148 N_C1_M1003_g N_Y_c_270_n 0.0102372f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_149 N_C1_c_179_n N_Y_c_274_n 9.1767e-19 $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_150 N_C1_c_177_n N_Y_c_274_n 0.0050009f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_151 N_C1_c_178_n N_Y_c_274_n 0.0159673f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_152 N_C1_c_179_n N_Y_c_275_n 0.0161324f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_153 N_C1_M1003_g N_VGND_c_338_n 0.00607661f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_154 N_C1_M1003_g N_VGND_c_343_n 0.00434272f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_155 N_C1_M1003_g N_VGND_c_344_n 0.00825192f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_156 N_VPWR_M1001_d N_A_156_368#_c_243_n 0.0087699f $X=1.23 $Y=1.84 $X2=0
+ $Y2=0
cc_157 N_VPWR_c_207_n N_A_156_368#_c_243_n 0.0297772f $X=1.47 $Y=2.76 $X2=0
+ $Y2=0
cc_158 N_VPWR_c_206_n N_A_156_368#_c_240_n 0.0469656f $X=0.48 $Y=2.455 $X2=0
+ $Y2=0
cc_159 N_VPWR_c_207_n N_A_156_368#_c_240_n 0.0139497f $X=1.47 $Y=2.76 $X2=0
+ $Y2=0
cc_160 N_VPWR_c_210_n N_A_156_368#_c_240_n 0.0145674f $X=1.265 $Y=3.33 $X2=0
+ $Y2=0
cc_161 N_VPWR_c_205_n N_A_156_368#_c_240_n 0.0119851f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_162 N_VPWR_c_207_n N_A_156_368#_c_241_n 0.0139497f $X=1.47 $Y=2.76 $X2=0
+ $Y2=0
cc_163 N_VPWR_c_212_n N_A_156_368#_c_241_n 0.0145674f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_164 N_VPWR_c_205_n N_A_156_368#_c_241_n 0.0119851f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_165 N_VPWR_M1001_d N_Y_c_286_n 0.0144403f $X=1.23 $Y=1.84 $X2=0 $Y2=0
cc_166 N_VPWR_c_212_n N_Y_c_275_n 0.0145938f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_167 N_VPWR_c_205_n N_Y_c_275_n 0.0120466f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_168 N_A_156_368#_M1000_d N_Y_c_286_n 0.00857291f $X=0.78 $Y=1.84 $X2=0 $Y2=0
cc_169 N_A_156_368#_M1007_d N_Y_c_286_n 0.0074438f $X=1.86 $Y=1.84 $X2=0 $Y2=0
cc_170 N_A_156_368#_c_243_n N_Y_c_286_n 0.0448167f $X=1.845 $Y=2.375 $X2=0 $Y2=0
cc_171 N_A_156_368#_c_240_n N_Y_c_286_n 0.0162525f $X=0.93 $Y=2.41 $X2=0 $Y2=0
cc_172 N_A_156_368#_c_241_n N_Y_c_286_n 0.0173542f $X=2.01 $Y=2.41 $X2=0 $Y2=0
cc_173 N_A_156_368#_c_240_n N_Y_c_281_n 0.00122866f $X=0.93 $Y=2.41 $X2=0 $Y2=0
cc_174 N_A_156_368#_c_241_n N_Y_c_275_n 0.0184959f $X=2.01 $Y=2.41 $X2=0 $Y2=0
cc_175 A_462_368# N_Y_c_286_n 0.010449f $X=2.31 $Y=1.84 $X2=2.775 $Y2=2.035
cc_176 N_Y_c_269_n N_VGND_M1009_d 0.00309832f $X=2.75 $Y=1.095 $X2=0 $Y2=0
cc_177 N_Y_c_272_n N_VGND_c_337_n 0.0189403f $X=2.04 $Y=0.765 $X2=0 $Y2=0
cc_178 N_Y_c_269_n N_VGND_c_338_n 0.024241f $X=2.75 $Y=1.095 $X2=0 $Y2=0
cc_179 N_Y_c_270_n N_VGND_c_338_n 0.0191903f $X=2.915 $Y=0.515 $X2=0 $Y2=0
cc_180 N_Y_c_272_n N_VGND_c_338_n 0.0196004f $X=2.04 $Y=0.765 $X2=0 $Y2=0
cc_181 N_Y_c_272_n N_VGND_c_341_n 0.0417862f $X=2.04 $Y=0.765 $X2=0 $Y2=0
cc_182 N_Y_c_270_n N_VGND_c_343_n 0.0145639f $X=2.915 $Y=0.515 $X2=0 $Y2=0
cc_183 N_Y_c_270_n N_VGND_c_344_n 0.0119984f $X=2.915 $Y=0.515 $X2=0 $Y2=0
cc_184 N_Y_c_272_n N_VGND_c_344_n 0.0341885f $X=2.04 $Y=0.765 $X2=0 $Y2=0
cc_185 N_Y_c_271_n A_159_74# 0.00366293f $X=1.085 $Y=0.765 $X2=-0.19 $Y2=-0.245
cc_186 N_Y_c_272_n A_231_74# 0.00122878f $X=2.04 $Y=0.765 $X2=-0.19 $Y2=-0.245
