# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__nor4bb_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__nor4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.180000 2.495000 1.540000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.265000 1.320000 1.315000 1.650000 ;
        RECT 1.085000 1.650000 1.315000 1.710000 ;
        RECT 1.085000 1.710000 2.890000 1.880000 ;
        RECT 2.720000 1.255000 3.920000 1.585000 ;
        RECT 2.720000 1.585000 2.890000 1.710000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.095000 1.530000 9.955000 1.860000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.125000 1.450000 10.455000 1.780000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.544200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.350000 0.945000 0.840000 ;
        RECT 0.615000 0.840000 2.915000 0.915000 ;
        RECT 0.615000 0.915000 5.775000 1.010000 ;
        RECT 0.615000 1.010000 0.945000 1.130000 ;
        RECT 1.615000 0.350000 1.945000 0.840000 ;
        RECT 2.665000 0.350000 2.915000 0.840000 ;
        RECT 2.665000 1.010000 5.775000 1.085000 ;
        RECT 3.595000 0.350000 3.845000 0.915000 ;
        RECT 4.515000 0.350000 4.845000 0.915000 ;
        RECT 5.525000 0.350000 5.775000 0.915000 ;
        RECT 5.525000 1.085000 5.775000 1.300000 ;
        RECT 5.525000 1.300000 6.615000 1.470000 ;
        RECT 5.990000 1.470000 6.320000 1.725000 ;
        RECT 5.990000 1.725000 7.230000 2.055000 ;
        RECT 6.445000 0.350000 6.775000 0.885000 ;
        RECT 6.445000 0.885000 8.035000 1.055000 ;
        RECT 6.445000 1.055000 6.615000 1.300000 ;
        RECT 7.705000 0.350000 8.035000 0.885000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  0.115000  0.085000  0.445000 1.130000 ;
        RECT  1.115000  0.085000  1.445000 0.670000 ;
        RECT  2.115000  0.085000  2.445000 0.670000 ;
        RECT  3.085000  0.085000  3.415000 0.745000 ;
        RECT  4.015000  0.085000  4.345000 0.745000 ;
        RECT  5.015000  0.085000  5.345000 0.745000 ;
        RECT  5.945000  0.085000  6.275000 1.130000 ;
        RECT  6.945000  0.085000  7.535000 0.680000 ;
        RECT  8.205000  0.085000  8.750000 0.680000 ;
        RECT 10.095000  0.085000 10.495000 0.940000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 11.040000 3.415000 ;
        RECT  1.115000 2.730000  1.445000 3.245000 ;
        RECT  2.065000 2.730000  2.435000 3.245000 ;
        RECT  8.790000 2.370000  9.120000 3.245000 ;
        RECT  9.775000 2.100000  9.945000 3.245000 ;
        RECT 10.595000 2.290000 10.925000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 1.820000  0.445000 2.050000 ;
      RECT  0.115000 2.050000  3.390000 2.220000 ;
      RECT  0.115000 2.220000  0.445000 2.980000 ;
      RECT  0.615000 2.390000  2.885000 2.560000 ;
      RECT  0.615000 2.560000  0.945000 2.980000 ;
      RECT  1.645000 2.560000  1.895000 2.980000 ;
      RECT  2.635000 2.560000  2.885000 2.905000 ;
      RECT  2.635000 2.905000  3.890000 3.075000 ;
      RECT  3.060000 1.755000  4.260000 1.925000 ;
      RECT  3.060000 1.925000  3.390000 2.050000 ;
      RECT  3.060000 2.220000  3.390000 2.735000 ;
      RECT  3.560000 2.095000  3.890000 2.905000 ;
      RECT  4.090000 1.925000  4.260000 2.905000 ;
      RECT  4.090000 2.905000  8.490000 3.075000 ;
      RECT  4.345000 1.255000  5.355000 1.585000 ;
      RECT  4.470000 1.755000  4.800000 2.565000 ;
      RECT  4.470000 2.565000  8.035000 2.735000 ;
      RECT  5.185000 1.585000  5.355000 2.225000 ;
      RECT  5.185000 2.225000  7.570000 2.395000 ;
      RECT  6.785000 1.225000  8.375000 1.555000 ;
      RECT  7.400000 1.725000  8.875000 1.895000 ;
      RECT  7.400000 1.895000  7.570000 2.225000 ;
      RECT  7.760000 2.065000  8.035000 2.565000 ;
      RECT  8.205000 0.850000  9.090000 1.020000 ;
      RECT  8.205000 1.020000  8.375000 1.225000 ;
      RECT  8.205000 2.065000  8.490000 2.905000 ;
      RECT  8.545000 1.190000  9.585000 1.360000 ;
      RECT  8.545000 1.360000  8.875000 1.725000 ;
      RECT  8.705000 1.895000  8.875000 2.030000 ;
      RECT  8.705000 2.030000  9.575000 2.200000 ;
      RECT  8.920000 0.255000  9.925000 0.425000 ;
      RECT  8.920000 0.425000  9.090000 0.850000 ;
      RECT  9.260000 0.670000  9.585000 1.190000 ;
      RECT  9.300000 2.200000  9.575000 2.980000 ;
      RECT  9.755000 0.425000  9.925000 1.110000 ;
      RECT  9.755000 1.110000 10.925000 1.280000 ;
      RECT 10.145000 1.950000 10.925000 2.120000 ;
      RECT 10.145000 2.120000 10.395000 2.980000 ;
      RECT 10.665000 0.350000 10.925000 1.110000 ;
      RECT 10.755000 1.280000 10.925000 1.950000 ;
  END
END sky130_fd_sc_hs__nor4bb_4
