* File: sky130_fd_sc_hs__a211o_1.spice
* Created: Tue Sep  1 19:48:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a211o_1.pex.spice"
.subckt sky130_fd_sc_hs__a211o_1  VNB VPB A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_81_264#_M1004_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.16776 AS=0.1961 PD=1.44783 PS=2.01 NRD=9.72 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1008 A_366_136# N_A2_M1008_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.64 AD=0.104
+ AS=0.14509 PD=0.965 PS=1.25217 NRD=20.148 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1009 N_A_81_264#_M1009_d N_A1_M1009_g A_366_136# VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.104 PD=0.92 PS=0.965 NRD=0 NRS=20.148 M=1 R=4.26667 SA=75001
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_B1_M1005_g N_A_81_264#_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1006 N_A_81_264#_M1006_d N_C1_M1006_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.112 PD=1.81 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75002
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_81_264#_M1000_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_279_392#_M1002_s VPB PSHORT L=0.15 W=1
+ AD=0.165 AS=0.275 PD=1.33 PS=2.55 NRD=4.9053 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1001 N_A_279_392#_M1001_d N_A1_M1001_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75000.7
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1003 A_550_392# N_B1_M1003_g N_A_279_392#_M1001_d VPB PSHORT L=0.15 W=1
+ AD=0.12 AS=0.15 PD=1.24 PS=1.3 NRD=12.7853 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1007 N_A_81_264#_M1007_d N_C1_M1007_g A_550_392# VPB PSHORT L=0.15 W=1
+ AD=0.275 AS=0.12 PD=2.55 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75001.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__a211o_1.pxi.spice"
*
.ends
*
*
