* NGSPICE file created from sky130_fd_sc_hs__nor2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor2b_2 A B_N VGND VNB VPB VPWR Y
M1000 Y a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.884e+11p pd=4.28e+06u as=7.744e+11p ps=6.56e+06u
M1001 Y a_27_392# a_228_368# VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=9.912e+11p ps=8.49e+06u
M1002 a_228_368# a_27_392# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A a_228_368# VPB pshort w=1.12e+06u l=150000u
+  ad=6.31e+11p pd=5.43e+06u as=0p ps=0u
M1004 a_228_368# A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1006 VGND a_27_392# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B_N a_27_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1008 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

