* File: sky130_fd_sc_hs__nand4b_2.pxi.spice
* Created: Thu Aug 27 20:52:14 2020
* 
x_PM_SKY130_FD_SC_HS__NAND4B_2%A_N N_A_N_M1015_g N_A_N_c_94_n N_A_N_c_98_n
+ N_A_N_M1003_g A_N A_N N_A_N_c_95_n N_A_N_c_96_n
+ PM_SKY130_FD_SC_HS__NAND4B_2%A_N
x_PM_SKY130_FD_SC_HS__NAND4B_2%A_27_74# N_A_27_74#_M1015_s N_A_27_74#_M1003_s
+ N_A_27_74#_c_134_n N_A_27_74#_M1009_g N_A_27_74#_M1008_g N_A_27_74#_c_135_n
+ N_A_27_74#_M1010_g N_A_27_74#_M1017_g N_A_27_74#_c_128_n N_A_27_74#_c_129_n
+ N_A_27_74#_c_130_n N_A_27_74#_c_136_n N_A_27_74#_c_137_n N_A_27_74#_c_138_n
+ N_A_27_74#_c_131_n N_A_27_74#_c_132_n N_A_27_74#_c_133_n
+ PM_SKY130_FD_SC_HS__NAND4B_2%A_27_74#
x_PM_SKY130_FD_SC_HS__NAND4B_2%B N_B_M1001_g N_B_c_216_n N_B_M1004_g N_B_M1014_g
+ N_B_c_217_n N_B_M1007_g B N_B_c_214_n N_B_c_215_n
+ PM_SKY130_FD_SC_HS__NAND4B_2%B
x_PM_SKY130_FD_SC_HS__NAND4B_2%C N_C_c_275_n N_C_M1002_g N_C_M1000_g N_C_c_276_n
+ N_C_M1005_g N_C_M1013_g C C N_C_c_274_n PM_SKY130_FD_SC_HS__NAND4B_2%C
x_PM_SKY130_FD_SC_HS__NAND4B_2%D N_D_c_332_n N_D_M1006_g N_D_M1011_g N_D_c_333_n
+ N_D_M1016_g N_D_M1012_g D D D N_D_c_331_n PM_SKY130_FD_SC_HS__NAND4B_2%D
x_PM_SKY130_FD_SC_HS__NAND4B_2%VPWR N_VPWR_M1003_d N_VPWR_M1010_s N_VPWR_M1007_s
+ N_VPWR_M1005_s N_VPWR_M1016_d N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_377_n
+ N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n
+ VPWR N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n
+ N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_374_n
+ PM_SKY130_FD_SC_HS__NAND4B_2%VPWR
x_PM_SKY130_FD_SC_HS__NAND4B_2%Y N_Y_M1008_s N_Y_M1009_d N_Y_M1004_d N_Y_M1002_d
+ N_Y_M1006_s N_Y_c_458_n N_Y_c_452_n N_Y_c_463_n N_Y_c_449_n N_Y_c_453_n
+ N_Y_c_494_n N_Y_c_454_n N_Y_c_499_n N_Y_c_514_n N_Y_c_455_n N_Y_c_450_n
+ N_Y_c_456_n N_Y_c_503_n Y Y PM_SKY130_FD_SC_HS__NAND4B_2%Y
x_PM_SKY130_FD_SC_HS__NAND4B_2%VGND N_VGND_M1015_d N_VGND_M1011_s N_VGND_c_551_n
+ N_VGND_c_552_n VGND N_VGND_c_553_n N_VGND_c_554_n N_VGND_c_555_n
+ N_VGND_c_556_n N_VGND_c_557_n N_VGND_c_558_n PM_SKY130_FD_SC_HS__NAND4B_2%VGND
x_PM_SKY130_FD_SC_HS__NAND4B_2%A_225_74# N_A_225_74#_M1008_d N_A_225_74#_M1017_d
+ N_A_225_74#_M1014_d N_A_225_74#_c_607_n N_A_225_74#_c_608_n
+ N_A_225_74#_c_609_n N_A_225_74#_c_621_n PM_SKY130_FD_SC_HS__NAND4B_2%A_225_74#
x_PM_SKY130_FD_SC_HS__NAND4B_2%A_490_74# N_A_490_74#_M1001_s N_A_490_74#_M1000_s
+ N_A_490_74#_c_644_n N_A_490_74#_c_650_n N_A_490_74#_c_645_n
+ PM_SKY130_FD_SC_HS__NAND4B_2%A_490_74#
x_PM_SKY130_FD_SC_HS__NAND4B_2%A_719_123# N_A_719_123#_M1000_d
+ N_A_719_123#_M1013_d N_A_719_123#_M1012_d N_A_719_123#_c_671_n
+ N_A_719_123#_c_672_n N_A_719_123#_c_673_n N_A_719_123#_c_674_n
+ N_A_719_123#_c_675_n N_A_719_123#_c_676_n N_A_719_123#_c_677_n
+ N_A_719_123#_c_678_n PM_SKY130_FD_SC_HS__NAND4B_2%A_719_123#
cc_1 VNB N_A_N_M1015_g 0.0318449f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_A_N_c_94_n 0.0132343f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.675
cc_3 VNB N_A_N_c_95_n 0.0245924f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_4 VNB N_A_N_c_96_n 0.0688411f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.345
cc_5 VNB N_A_27_74#_M1008_g 0.0266096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_74#_M1017_g 0.0239157f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.345
cc_7 VNB N_A_27_74#_c_128_n 0.0203664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_129_n 0.0105263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_130_n 0.00949248f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_10 VNB N_A_27_74#_c_131_n 0.00567489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_132_n 0.00646829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_133_n 0.0381438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_M1001_g 0.0255964f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_14 VNB N_B_M1014_g 0.0293822f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_B_c_214_n 0.00465678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_215_n 0.0553056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_M1000_g 0.023676f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.675
cc_18 VNB N_C_M1013_g 0.0200129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB C 0.00377768f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_20 VNB N_C_c_274_n 0.0573263f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.345
cc_21 VNB N_D_M1011_g 0.0202431f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.675
cc_22 VNB N_D_M1012_g 0.028245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB D 0.0203907f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_24 VNB N_D_c_331_n 0.036671f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_25 VNB N_VPWR_c_374_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_449_n 0.00841801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_450_n 0.00418682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 0.0025475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_551_n 0.0100536f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.34
cc_30 VNB N_VGND_c_552_n 0.0069637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_553_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_32 VNB N_VGND_c_554_n 0.0979637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_555_n 0.0183664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_556_n 0.332581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_557_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_558_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_225_74#_c_607_n 0.00846754f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_38 VNB N_A_225_74#_c_608_n 0.00194367f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_39 VNB N_A_225_74#_c_609_n 0.00305483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_490_74#_c_644_n 0.0219302f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.765
cc_41 VNB N_A_490_74#_c_645_n 0.00366476f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_42 VNB N_A_719_123#_c_671_n 0.00392221f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_43 VNB N_A_719_123#_c_672_n 0.00551296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_719_123#_c_673_n 0.00461713f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.345
cc_45 VNB N_A_719_123#_c_674_n 0.00210056f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_46 VNB N_A_719_123#_c_675_n 0.00326619f $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=1.345
cc_47 VNB N_A_719_123#_c_676_n 0.0131055f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.345
cc_48 VNB N_A_719_123#_c_677_n 0.0220272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_719_123#_c_678_n 0.00178419f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_50 VPB N_A_N_c_94_n 0.00124349f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.675
cc_51 VPB N_A_N_c_98_n 0.0261592f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.765
cc_52 VPB N_A_27_74#_c_134_n 0.017213f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.765
cc_53 VPB N_A_27_74#_c_135_n 0.0179154f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.345
cc_54 VPB N_A_27_74#_c_136_n 0.0416815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_74#_c_137_n 0.00256945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_74#_c_138_n 0.0094432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_74#_c_132_n 0.00467504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_27_74#_c_133_n 0.0231746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_B_c_216_n 0.0178086f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.51
cc_60 VPB N_B_c_217_n 0.0157968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_B_c_214_n 0.00720788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B_c_215_n 0.0312883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_C_c_275_n 0.0164756f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.18
cc_64 VPB N_C_c_276_n 0.0171347f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=2.34
cc_65 VPB C 0.00496447f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.345
cc_66 VPB N_C_c_274_n 0.0231586f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.345
cc_67 VPB N_D_c_332_n 0.0170595f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.18
cc_68 VPB N_D_c_333_n 0.0179656f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=2.34
cc_69 VPB D 0.0159088f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.345
cc_70 VPB N_D_c_331_n 0.0210926f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.345
cc_71 VPB N_VPWR_c_375_n 0.0104692f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.345
cc_72 VPB N_VPWR_c_376_n 0.0110056f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.345
cc_73 VPB N_VPWR_c_377_n 0.00900305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_378_n 0.00988376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_379_n 0.0113253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_380_n 0.0508411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_381_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_382_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_383_n 0.0332141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_384_n 0.0175344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_385_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_386_n 0.0199677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_387_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_388_n 0.0114188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_389_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_374_n 0.0943814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_Y_c_452_n 0.00239217f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.345
cc_88 VPB N_Y_c_453_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.345
cc_89 VPB N_Y_c_454_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_Y_c_455_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_Y_c_456_n 0.00223019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB Y 0.00184384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 N_A_N_c_98_n N_A_27_74#_c_134_n 0.01564f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_N_c_96_n N_A_27_74#_M1008_g 0.00377133f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_95 N_A_N_M1015_g N_A_27_74#_c_128_n 0.00264672f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_96 N_A_N_M1015_g N_A_27_74#_c_129_n 0.0143914f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_97 N_A_N_c_95_n N_A_27_74#_c_129_n 0.0415659f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_98 N_A_N_c_96_n N_A_27_74#_c_129_n 0.00985512f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_99 N_A_N_c_95_n N_A_27_74#_c_130_n 0.0204809f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_100 N_A_N_c_96_n N_A_27_74#_c_130_n 0.00115581f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_101 N_A_N_c_98_n N_A_27_74#_c_136_n 0.0125615f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_N_c_98_n N_A_27_74#_c_137_n 0.012624f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A_N_c_95_n N_A_27_74#_c_137_n 0.010678f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_104 N_A_N_c_98_n N_A_27_74#_c_138_n 0.00436428f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_N_c_95_n N_A_27_74#_c_138_n 0.0276947f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_106 N_A_N_c_96_n N_A_27_74#_c_138_n 0.00724507f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_107 N_A_N_M1015_g N_A_27_74#_c_131_n 0.0037584f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_108 N_A_N_c_95_n N_A_27_74#_c_131_n 0.013468f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_109 N_A_N_c_96_n N_A_27_74#_c_131_n 5.96187e-19 $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_110 N_A_N_c_95_n N_A_27_74#_c_132_n 0.013971f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_111 N_A_N_c_96_n N_A_27_74#_c_132_n 0.00529557f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_112 N_A_N_c_96_n N_A_27_74#_c_133_n 0.0126129f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_113 N_A_N_c_98_n N_VPWR_c_375_n 0.0107596f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_N_c_98_n N_VPWR_c_383_n 0.00481995f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_N_c_98_n N_VPWR_c_374_n 0.00508379f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_N_M1015_g N_VGND_c_551_n 0.0115915f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_117 N_A_N_M1015_g N_VGND_c_553_n 0.00383152f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_118 N_A_N_M1015_g N_VGND_c_556_n 0.00387625f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_119 N_A_N_M1015_g N_A_225_74#_c_607_n 6.17645e-19 $X=0.495 $Y=0.69 $X2=0
+ $Y2=0
cc_120 N_A_27_74#_M1017_g N_B_M1001_g 0.0334156f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_27_74#_c_135_n N_B_c_216_n 0.0102632f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_27_74#_c_135_n N_B_c_214_n 4.53592e-19 $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_27_74#_c_132_n N_B_c_214_n 0.017469f $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_27_74#_c_133_n N_B_c_214_n 0.0069357f $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_125 N_A_27_74#_c_132_n N_B_c_215_n 2.0756e-19 $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A_27_74#_c_133_n N_B_c_215_n 0.0189662f $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_127 N_A_27_74#_c_137_n N_VPWR_M1003_d 0.00173539f $X=1.155 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_27_74#_c_132_n N_VPWR_M1003_d 0.0016378f $X=1.555 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_27_74#_c_134_n N_VPWR_c_375_n 0.0138446f $X=1.435 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_27_74#_c_135_n N_VPWR_c_375_n 6.08654e-19 $X=1.885 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_27_74#_c_136_n N_VPWR_c_375_n 0.0564881f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_27_74#_c_137_n N_VPWR_c_375_n 0.0092384f $X=1.155 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_27_74#_c_132_n N_VPWR_c_375_n 0.014575f $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A_27_74#_c_135_n N_VPWR_c_376_n 0.00248287f $X=1.885 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_27_74#_c_136_n N_VPWR_c_383_n 0.0097982f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_27_74#_c_134_n N_VPWR_c_384_n 0.00429299f $X=1.435 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_27_74#_c_135_n N_VPWR_c_384_n 0.00445602f $X=1.885 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_27_74#_c_134_n N_VPWR_c_374_n 0.00847721f $X=1.435 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_27_74#_c_135_n N_VPWR_c_374_n 0.00859404f $X=1.885 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_27_74#_c_136_n N_VPWR_c_374_n 0.0111907f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_27_74#_c_135_n N_Y_c_458_n 0.00479881f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_27_74#_c_132_n N_Y_c_458_n 0.0133428f $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A_27_74#_c_133_n N_Y_c_458_n 0.00318959f $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_144 N_A_27_74#_c_134_n N_Y_c_452_n 2.48635e-19 $X=1.435 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_27_74#_c_135_n N_Y_c_452_n 0.0144534f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_27_74#_c_135_n N_Y_c_463_n 0.0173717f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_27_74#_c_133_n N_Y_c_463_n 0.00102375f $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_148 N_A_27_74#_M1017_g N_Y_c_449_n 0.0129671f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_27_74#_M1008_g N_Y_c_450_n 0.00727448f $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_27_74#_M1017_g N_Y_c_450_n 0.00682377f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_27_74#_c_129_n N_Y_c_450_n 0.0119985f $X=1.155 $Y=0.925 $X2=0 $Y2=0
cc_152 N_A_27_74#_c_131_n N_Y_c_450_n 0.0108039f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_153 N_A_27_74#_c_132_n N_Y_c_450_n 0.0147728f $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A_27_74#_c_133_n N_Y_c_450_n 0.00225444f $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_155 N_A_27_74#_c_129_n N_VGND_M1015_d 0.00425898f $X=1.155 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_27_74#_M1008_g N_VGND_c_551_n 0.0032818f $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_27_74#_c_128_n N_VGND_c_551_n 0.0121972f $X=0.28 $Y=0.68 $X2=0 $Y2=0
cc_158 N_A_27_74#_c_129_n N_VGND_c_551_n 0.0215034f $X=1.155 $Y=0.925 $X2=0
+ $Y2=0
cc_159 N_A_27_74#_c_128_n N_VGND_c_553_n 0.0110419f $X=0.28 $Y=0.68 $X2=0 $Y2=0
cc_160 N_A_27_74#_M1008_g N_VGND_c_554_n 0.00291649f $X=1.485 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_27_74#_M1017_g N_VGND_c_554_n 0.00291649f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_162 N_A_27_74#_M1008_g N_VGND_c_556_n 0.00364413f $X=1.485 $Y=0.74 $X2=0
+ $Y2=0
cc_163 N_A_27_74#_M1017_g N_VGND_c_556_n 0.00359511f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_164 N_A_27_74#_c_128_n N_VGND_c_556_n 0.00915013f $X=0.28 $Y=0.68 $X2=0 $Y2=0
cc_165 N_A_27_74#_c_129_n N_VGND_c_556_n 0.0144197f $X=1.155 $Y=0.925 $X2=0
+ $Y2=0
cc_166 N_A_27_74#_c_129_n N_A_225_74#_M1008_d 0.00509711f $X=1.155 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_167 N_A_27_74#_c_131_n N_A_225_74#_M1008_d 0.00174945f $X=1.24 $Y=1.35
+ $X2=-0.19 $Y2=-0.245
cc_168 N_A_27_74#_M1008_g N_A_225_74#_c_607_n 0.0154696f $X=1.485 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_27_74#_M1017_g N_A_225_74#_c_607_n 0.0122685f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_27_74#_c_129_n N_A_225_74#_c_607_n 0.0148275f $X=1.155 $Y=0.925 $X2=0
+ $Y2=0
cc_171 N_B_c_217_n N_C_c_275_n 0.0304769f $X=3.15 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_172 N_B_c_215_n C 0.00326268f $X=2.965 $Y=1.557 $X2=0 $Y2=0
cc_173 N_B_c_215_n N_C_c_274_n 0.0174382f $X=2.965 $Y=1.557 $X2=0 $Y2=0
cc_174 N_B_c_216_n N_VPWR_c_376_n 0.00254884f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_175 N_B_c_217_n N_VPWR_c_377_n 0.00598632f $X=3.15 $Y=1.765 $X2=0 $Y2=0
cc_176 N_B_c_216_n N_VPWR_c_381_n 0.00445602f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_177 N_B_c_217_n N_VPWR_c_381_n 0.00445602f $X=3.15 $Y=1.765 $X2=0 $Y2=0
cc_178 N_B_c_216_n N_VPWR_c_374_n 0.00859404f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_179 N_B_c_217_n N_VPWR_c_374_n 0.00857825f $X=3.15 $Y=1.765 $X2=0 $Y2=0
cc_180 N_B_c_216_n N_Y_c_463_n 0.0177366f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_181 N_B_c_214_n N_Y_c_463_n 0.0426108f $X=2.425 $Y=1.515 $X2=0 $Y2=0
cc_182 N_B_c_215_n N_Y_c_463_n 0.00174282f $X=2.965 $Y=1.557 $X2=0 $Y2=0
cc_183 N_B_M1001_g N_Y_c_449_n 0.0112328f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_184 N_B_M1014_g N_Y_c_449_n 0.0132383f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_185 N_B_c_214_n N_Y_c_449_n 0.042165f $X=2.425 $Y=1.515 $X2=0 $Y2=0
cc_186 N_B_c_215_n N_Y_c_449_n 0.0101219f $X=2.965 $Y=1.557 $X2=0 $Y2=0
cc_187 N_B_c_216_n N_Y_c_453_n 0.0150799f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_188 N_B_c_217_n N_Y_c_453_n 0.0109514f $X=3.15 $Y=1.765 $X2=0 $Y2=0
cc_189 N_B_c_217_n N_Y_c_454_n 6.63528e-19 $X=3.15 $Y=1.765 $X2=0 $Y2=0
cc_190 N_B_M1001_g N_Y_c_450_n 9.39477e-19 $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_191 N_B_c_216_n N_Y_c_456_n 0.00713046f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_192 N_B_c_217_n N_Y_c_456_n 0.0131453f $X=3.15 $Y=1.765 $X2=0 $Y2=0
cc_193 N_B_c_215_n N_Y_c_456_n 0.00805211f $X=2.965 $Y=1.557 $X2=0 $Y2=0
cc_194 N_B_M1001_g Y 7.76767e-19 $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_195 N_B_c_216_n Y 9.32952e-19 $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_196 N_B_M1014_g Y 0.00655125f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_197 N_B_c_217_n Y 0.00134606f $X=3.15 $Y=1.765 $X2=0 $Y2=0
cc_198 N_B_c_214_n Y 0.0166917f $X=2.425 $Y=1.515 $X2=0 $Y2=0
cc_199 N_B_c_215_n Y 0.0255068f $X=2.965 $Y=1.557 $X2=0 $Y2=0
cc_200 N_B_M1001_g N_VGND_c_554_n 0.00324657f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_201 N_B_M1014_g N_VGND_c_554_n 0.00278271f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B_M1001_g N_VGND_c_556_n 0.00412223f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_203 N_B_M1014_g N_VGND_c_556_n 0.00359811f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_204 N_B_M1001_g N_A_225_74#_c_608_n 0.00739353f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B_M1014_g N_A_225_74#_c_608_n 9.2292e-19 $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B_M1001_g N_A_225_74#_c_609_n 3.34639e-19 $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B_M1014_g N_A_225_74#_c_609_n 0.00257863f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B_c_215_n N_A_225_74#_c_609_n 7.58336e-19 $X=2.965 $Y=1.557 $X2=0 $Y2=0
cc_209 N_B_M1001_g N_A_225_74#_c_621_n 0.00982687f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B_M1014_g N_A_225_74#_c_621_n 0.00850118f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B_M1014_g N_A_490_74#_c_644_n 0.0120769f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B_M1001_g N_A_490_74#_c_645_n 0.00416113f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B_M1014_g N_A_719_123#_c_671_n 0.00139553f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B_M1014_g N_A_719_123#_c_673_n 0.00312109f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_215 N_C_c_276_n N_D_c_332_n 0.0237503f $X=4.15 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_216 N_C_M1013_g N_D_M1011_g 0.011802f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_217 C D 0.0279008f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_218 N_C_c_274_n D 0.0079955f $X=4.15 $Y=1.557 $X2=0 $Y2=0
cc_219 C N_D_c_331_n 3.13064e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_220 N_C_c_274_n N_D_c_331_n 0.0168681f $X=4.15 $Y=1.557 $X2=0 $Y2=0
cc_221 N_C_c_275_n N_VPWR_c_377_n 0.00737447f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_222 N_C_c_276_n N_VPWR_c_378_n 0.0101544f $X=4.15 $Y=1.765 $X2=0 $Y2=0
cc_223 N_C_c_275_n N_VPWR_c_385_n 0.00445602f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_224 N_C_c_276_n N_VPWR_c_385_n 0.00445602f $X=4.15 $Y=1.765 $X2=0 $Y2=0
cc_225 N_C_c_275_n N_VPWR_c_374_n 0.00857825f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_226 N_C_c_276_n N_VPWR_c_374_n 0.00859856f $X=4.15 $Y=1.765 $X2=0 $Y2=0
cc_227 N_C_M1000_g N_Y_c_449_n 5.99596e-19 $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_228 N_C_c_275_n N_Y_c_453_n 6.63528e-19 $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_229 N_C_c_275_n N_Y_c_494_n 0.012262f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_230 C N_Y_c_494_n 0.0188972f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_231 N_C_c_274_n N_Y_c_494_n 3.87644e-19 $X=4.15 $Y=1.557 $X2=0 $Y2=0
cc_232 N_C_c_275_n N_Y_c_454_n 0.0104413f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_233 N_C_c_276_n N_Y_c_454_n 0.0117453f $X=4.15 $Y=1.765 $X2=0 $Y2=0
cc_234 N_C_c_276_n N_Y_c_499_n 0.0137046f $X=4.15 $Y=1.765 $X2=0 $Y2=0
cc_235 C N_Y_c_499_n 0.00762725f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_236 N_C_c_274_n N_Y_c_499_n 0.00584887f $X=4.15 $Y=1.557 $X2=0 $Y2=0
cc_237 N_C_c_276_n N_Y_c_455_n 8.65319e-19 $X=4.15 $Y=1.765 $X2=0 $Y2=0
cc_238 N_C_c_275_n N_Y_c_503_n 4.27055e-19 $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_239 N_C_c_276_n N_Y_c_503_n 4.27055e-19 $X=4.15 $Y=1.765 $X2=0 $Y2=0
cc_240 C N_Y_c_503_n 0.0237598f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_241 N_C_c_274_n N_Y_c_503_n 0.00144091f $X=4.15 $Y=1.557 $X2=0 $Y2=0
cc_242 N_C_c_275_n Y 0.00148392f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_243 N_C_M1000_g Y 0.00367138f $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_244 C Y 0.0265881f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_245 N_C_c_274_n Y 4.81621e-19 $X=4.15 $Y=1.557 $X2=0 $Y2=0
cc_246 N_C_M1013_g N_VGND_c_552_n 4.25532e-19 $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_247 N_C_M1000_g N_VGND_c_554_n 8.94875e-19 $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_248 N_C_M1013_g N_VGND_c_554_n 0.00465842f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_249 N_C_M1013_g N_VGND_c_556_n 0.00441603f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_250 N_C_M1000_g N_A_490_74#_c_644_n 0.011917f $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_251 N_C_M1013_g N_A_490_74#_c_644_n 0.00409781f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_252 N_C_M1000_g N_A_490_74#_c_650_n 0.00944526f $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_253 N_C_M1013_g N_A_490_74#_c_650_n 0.00370415f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_254 N_C_M1000_g N_A_719_123#_c_672_n 0.0140147f $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_255 N_C_M1013_g N_A_719_123#_c_672_n 0.0183977f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_256 C N_A_719_123#_c_672_n 0.0285914f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_257 N_C_c_274_n N_A_719_123#_c_672_n 0.0043122f $X=4.15 $Y=1.557 $X2=0 $Y2=0
cc_258 C N_A_719_123#_c_673_n 0.0212141f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_259 N_C_c_274_n N_A_719_123#_c_673_n 0.00641319f $X=4.15 $Y=1.557 $X2=0 $Y2=0
cc_260 N_C_M1013_g N_A_719_123#_c_674_n 3.98786e-19 $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_261 N_D_c_332_n N_VPWR_c_378_n 0.0103027f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_262 N_D_c_333_n N_VPWR_c_380_n 0.00506392f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_263 D N_VPWR_c_380_n 0.0232961f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_264 N_D_c_332_n N_VPWR_c_386_n 0.00445602f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_265 N_D_c_333_n N_VPWR_c_386_n 0.00445602f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_266 N_D_c_332_n N_VPWR_c_374_n 0.00859408f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_267 N_D_c_333_n N_VPWR_c_374_n 0.00860428f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_268 N_D_c_332_n N_Y_c_454_n 8.77392e-19 $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_269 N_D_c_332_n N_Y_c_499_n 0.0128325f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_270 D N_Y_c_499_n 0.0300484f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_271 N_D_c_332_n N_Y_c_514_n 4.27055e-19 $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_272 N_D_c_333_n N_Y_c_514_n 0.0019041f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_273 D N_Y_c_514_n 0.0237598f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_274 N_D_c_331_n N_Y_c_514_n 0.00144303f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_275 N_D_c_332_n N_Y_c_455_n 0.0114079f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_276 N_D_c_333_n N_Y_c_455_n 0.00906641f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_277 N_D_M1011_g N_VGND_c_552_n 0.00804216f $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_278 N_D_M1012_g N_VGND_c_552_n 0.00985076f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_279 N_D_M1011_g N_VGND_c_554_n 0.00449979f $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_280 N_D_M1012_g N_VGND_c_555_n 0.00522181f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_281 N_D_M1011_g N_VGND_c_556_n 0.00445136f $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_282 N_D_M1012_g N_VGND_c_556_n 0.00515793f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_283 N_D_M1011_g N_A_490_74#_c_644_n 3.29564e-19 $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_284 D N_A_719_123#_c_672_n 0.00483207f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_285 N_D_M1011_g N_A_719_123#_c_674_n 3.99083e-19 $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_286 N_D_M1011_g N_A_719_123#_c_675_n 0.0148218f $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_287 N_D_M1012_g N_A_719_123#_c_675_n 0.0154779f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_288 D N_A_719_123#_c_675_n 0.0544516f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_289 N_D_c_331_n N_A_719_123#_c_675_n 0.002768f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_290 D N_A_719_123#_c_676_n 0.0216404f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_291 N_D_M1012_g N_A_719_123#_c_677_n 0.0015993f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_292 D N_A_719_123#_c_678_n 0.017132f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_293 N_VPWR_c_375_n N_Y_c_452_n 0.0315621f $X=1.205 $Y=2.105 $X2=0 $Y2=0
cc_294 N_VPWR_c_376_n N_Y_c_452_n 0.0260414f $X=2.475 $Y=2.455 $X2=0 $Y2=0
cc_295 N_VPWR_c_384_n N_Y_c_452_n 0.0121397f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_c_374_n N_Y_c_452_n 0.0100153f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_297 N_VPWR_M1010_s N_Y_c_463_n 0.014615f $X=1.96 $Y=1.84 $X2=0 $Y2=0
cc_298 N_VPWR_c_376_n N_Y_c_463_n 0.0448286f $X=2.475 $Y=2.455 $X2=0 $Y2=0
cc_299 N_VPWR_c_376_n N_Y_c_453_n 0.0267545f $X=2.475 $Y=2.455 $X2=0 $Y2=0
cc_300 N_VPWR_c_377_n N_Y_c_453_n 0.0266809f $X=3.425 $Y=2.415 $X2=0 $Y2=0
cc_301 N_VPWR_c_381_n N_Y_c_453_n 0.014552f $X=3.26 $Y=3.33 $X2=0 $Y2=0
cc_302 N_VPWR_c_374_n N_Y_c_453_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_303 N_VPWR_M1007_s N_Y_c_494_n 0.0119577f $X=3.225 $Y=1.84 $X2=0 $Y2=0
cc_304 N_VPWR_c_377_n N_Y_c_494_n 0.0232685f $X=3.425 $Y=2.415 $X2=0 $Y2=0
cc_305 N_VPWR_c_377_n N_Y_c_454_n 0.0266809f $X=3.425 $Y=2.415 $X2=0 $Y2=0
cc_306 N_VPWR_c_378_n N_Y_c_454_n 0.0424981f $X=4.485 $Y=2.41 $X2=0 $Y2=0
cc_307 N_VPWR_c_385_n N_Y_c_454_n 0.014552f $X=4.32 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_374_n N_Y_c_454_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_M1005_s N_Y_c_499_n 0.0117594f $X=4.225 $Y=1.84 $X2=0 $Y2=0
cc_310 N_VPWR_c_378_n N_Y_c_499_n 0.0266856f $X=4.485 $Y=2.41 $X2=0 $Y2=0
cc_311 N_VPWR_c_378_n N_Y_c_455_n 0.0455583f $X=4.485 $Y=2.41 $X2=0 $Y2=0
cc_312 N_VPWR_c_380_n N_Y_c_455_n 0.0330049f $X=5.475 $Y=2.115 $X2=0 $Y2=0
cc_313 N_VPWR_c_386_n N_Y_c_455_n 0.014552f $X=5.36 $Y=3.33 $X2=0 $Y2=0
cc_314 N_VPWR_c_374_n N_Y_c_455_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_315 N_Y_c_449_n N_A_225_74#_M1017_d 0.00176461f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_316 N_Y_c_449_n N_A_225_74#_M1014_d 0.00300606f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_317 N_Y_M1008_s N_A_225_74#_c_607_n 0.00211578f $X=1.56 $Y=0.37 $X2=0 $Y2=0
cc_318 N_Y_c_449_n N_A_225_74#_c_607_n 0.00459468f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_319 N_Y_c_450_n N_A_225_74#_c_607_n 0.0187497f $X=1.715 $Y=0.965 $X2=0 $Y2=0
cc_320 N_Y_c_449_n N_A_225_74#_c_608_n 0.0149311f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_321 N_Y_c_449_n N_A_225_74#_c_621_n 0.0540678f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_322 N_Y_c_449_n N_A_490_74#_M1001_s 0.00391227f $X=3.005 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_323 N_Y_c_449_n N_A_719_123#_c_673_n 0.00962672f $X=3.005 $Y=1.095 $X2=0
+ $Y2=0
cc_324 N_VGND_c_551_n N_A_225_74#_c_607_n 0.0198879f $X=0.71 $Y=0.55 $X2=0 $Y2=0
cc_325 N_VGND_c_554_n N_A_225_74#_c_607_n 0.039681f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_556_n N_A_225_74#_c_607_n 0.0333579f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_554_n N_A_225_74#_c_608_n 0.0107387f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_556_n N_A_225_74#_c_608_n 0.00894442f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_329 N_VGND_c_554_n N_A_225_74#_c_621_n 0.00237563f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_330 N_VGND_c_556_n N_A_225_74#_c_621_n 0.00539332f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_331 N_VGND_c_552_n N_A_490_74#_c_644_n 0.00485382f $X=5.03 $Y=0.58 $X2=0
+ $Y2=0
cc_332 N_VGND_c_554_n N_A_490_74#_c_644_n 0.0231371f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_556_n N_A_490_74#_c_644_n 0.0127322f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_334 N_VGND_c_554_n N_A_490_74#_c_645_n 0.0966814f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_335 N_VGND_c_556_n N_A_490_74#_c_645_n 0.0558053f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_336 N_VGND_c_552_n N_A_719_123#_c_674_n 0.0142351f $X=5.03 $Y=0.58 $X2=0
+ $Y2=0
cc_337 N_VGND_c_554_n N_A_719_123#_c_674_n 0.00698151f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_338 N_VGND_c_556_n N_A_719_123#_c_674_n 0.00673015f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_M1011_s N_A_719_123#_c_675_n 0.00200085f $X=4.89 $Y=0.42 $X2=0
+ $Y2=0
cc_340 N_VGND_c_552_n N_A_719_123#_c_675_n 0.017643f $X=5.03 $Y=0.58 $X2=0 $Y2=0
cc_341 N_VGND_c_552_n N_A_719_123#_c_677_n 0.0125364f $X=5.03 $Y=0.58 $X2=0
+ $Y2=0
cc_342 N_VGND_c_555_n N_A_719_123#_c_677_n 0.00920966f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_343 N_VGND_c_556_n N_A_719_123#_c_677_n 0.00887807f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_344 N_A_225_74#_c_621_n N_A_490_74#_M1001_s 0.00727678f $X=3.015 $Y=0.717
+ $X2=-0.19 $Y2=-0.245
cc_345 N_A_225_74#_M1014_d N_A_490_74#_c_644_n 0.00226585f $X=3.04 $Y=0.37 $X2=0
+ $Y2=0
cc_346 N_A_225_74#_c_609_n N_A_490_74#_c_644_n 0.0191024f $X=3.18 $Y=0.715 $X2=0
+ $Y2=0
cc_347 N_A_225_74#_c_621_n N_A_490_74#_c_644_n 0.00570513f $X=3.015 $Y=0.717
+ $X2=0 $Y2=0
cc_348 N_A_225_74#_c_608_n N_A_490_74#_c_645_n 0.00599132f $X=2.2 $Y=0.49 $X2=0
+ $Y2=0
cc_349 N_A_225_74#_c_621_n N_A_490_74#_c_645_n 0.0232532f $X=3.015 $Y=0.717
+ $X2=0 $Y2=0
cc_350 N_A_225_74#_c_609_n N_A_719_123#_c_671_n 0.0167582f $X=3.18 $Y=0.715
+ $X2=0 $Y2=0
cc_351 N_A_490_74#_c_644_n N_A_719_123#_M1000_d 0.00206713f $X=4.005 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_352 N_A_490_74#_c_644_n N_A_719_123#_c_671_n 0.0187376f $X=4.005 $Y=0.34
+ $X2=0 $Y2=0
cc_353 N_A_490_74#_M1000_s N_A_719_123#_c_672_n 0.00178571f $X=4.03 $Y=0.42
+ $X2=0 $Y2=0
cc_354 N_A_490_74#_c_644_n N_A_719_123#_c_672_n 0.00356278f $X=4.005 $Y=0.34
+ $X2=0 $Y2=0
cc_355 N_A_490_74#_c_650_n N_A_719_123#_c_672_n 0.0171301f $X=4.17 $Y=0.58 $X2=0
+ $Y2=0
cc_356 N_A_490_74#_c_644_n N_A_719_123#_c_674_n 0.00178319f $X=4.005 $Y=0.34
+ $X2=0 $Y2=0
