* File: sky130_fd_sc_hs__o22ai_2.pex.spice
* Created: Thu Aug 27 21:00:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O22AI_2%B1 3 5 7 8 10 13 15 16 17 26
c46 17 0 1.08831e-19 $X=1.2 $Y=1.665
c47 8 0 1.00781e-20 $X=1.01 $Y=1.765
c48 5 0 9.04372e-20 $X=0.51 $Y=1.765
r49 26 27 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=1.01 $Y=1.557
+ $X2=1.025 $Y2=1.557
r50 24 26 10.9253 $w=3.75e-07 $l=8.5e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=1.01 $Y2=1.557
r51 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.515 $X2=0.925 $Y2=1.515
r52 22 24 53.3413 $w=3.75e-07 $l=4.15e-07 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.925 $Y2=1.557
r53 21 22 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r54 17 25 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.925 $Y2=1.565
r55 16 25 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.925 $Y2=1.565
r56 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r57 11 27 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.025 $Y=1.35
+ $X2=1.025 $Y2=1.557
r58 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.025 $Y=1.35
+ $X2=1.025 $Y2=0.74
r59 8 26 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.01 $Y=1.765
+ $X2=1.01 $Y2=1.557
r60 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.01 $Y=1.765
+ $X2=1.01 $Y2=2.4
r61 5 22 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r62 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r63 1 21 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r64 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%B2 1 3 6 8 10 13 15 21 22
c57 21 0 1.00781e-20 $X=1.65 $Y=1.515
c58 13 0 1.81856e-19 $X=1.995 $Y=0.74
c59 1 0 1.08831e-19 $X=1.46 $Y=1.765
r60 22 23 11.5408 $w=3.55e-07 $l=8.5e-08 $layer=POLY_cond $X=1.91 $Y=1.557
+ $X2=1.995 $Y2=1.557
r61 20 22 35.3014 $w=3.55e-07 $l=2.6e-07 $layer=POLY_cond $X=1.65 $Y=1.557
+ $X2=1.91 $Y2=1.557
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r63 18 20 21.0451 $w=3.55e-07 $l=1.55e-07 $layer=POLY_cond $X=1.495 $Y=1.557
+ $X2=1.65 $Y2=1.557
r64 17 18 4.75211 $w=3.55e-07 $l=3.5e-08 $layer=POLY_cond $X=1.46 $Y=1.557
+ $X2=1.495 $Y2=1.557
r65 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.515
r66 11 23 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.995 $Y=1.35
+ $X2=1.995 $Y2=1.557
r67 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.995 $Y=1.35
+ $X2=1.995 $Y2=0.74
r68 8 22 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=1.557
r69 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=2.4
r70 4 18 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=1.557
r71 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=0.74
r72 1 17 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.46 $Y2=1.557
r73 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.46 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%A2 3 5 7 8 10 13 17 23 24
c61 23 0 1.81856e-19 $X=3.17 $Y=1.465
c62 17 0 1.37374e-19 $X=3.6 $Y=1.665
c63 8 0 1.88367e-19 $X=3.37 $Y=1.765
r64 24 25 0.616368 $w=3.91e-07 $l=5e-09 $layer=POLY_cond $X=3.37 $Y=1.532
+ $X2=3.375 $Y2=1.532
r65 22 24 24.6547 $w=3.91e-07 $l=2e-07 $layer=POLY_cond $X=3.17 $Y=1.532
+ $X2=3.37 $Y2=1.532
r66 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.17
+ $Y=1.465 $X2=3.17 $Y2=1.465
r67 20 22 30.8184 $w=3.91e-07 $l=2.5e-07 $layer=POLY_cond $X=2.92 $Y=1.532
+ $X2=3.17 $Y2=1.532
r68 19 20 1.8491 $w=3.91e-07 $l=1.5e-08 $layer=POLY_cond $X=2.905 $Y=1.532
+ $X2=2.92 $Y2=1.532
r69 17 23 15.897 $w=3.3e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.54 $X2=3.17
+ $Y2=1.54
r70 11 25 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.375 $Y=1.3
+ $X2=3.375 $Y2=1.532
r71 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.375 $Y=1.3
+ $X2=3.375 $Y2=0.74
r72 8 24 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.37 $Y=1.765
+ $X2=3.37 $Y2=1.532
r73 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.37 $Y=1.765
+ $X2=3.37 $Y2=2.4
r74 5 20 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.92 $Y=1.765
+ $X2=2.92 $Y2=1.532
r75 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.92 $Y=1.765
+ $X2=2.92 $Y2=2.4
r76 1 19 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.905 $Y=1.3
+ $X2=2.905 $Y2=1.532
r77 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.905 $Y=1.3 $X2=2.905
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%A1 3 5 7 8 10 13 15 16 22
c47 5 0 1.37374e-19 $X=3.82 $Y=1.765
r48 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.415
+ $Y=1.515 $X2=4.415 $Y2=1.515
r49 22 24 14.4863 $w=3.66e-07 $l=1.1e-07 $layer=POLY_cond $X=4.305 $Y=1.557
+ $X2=4.415 $Y2=1.557
r50 21 22 4.60929 $w=3.66e-07 $l=3.5e-08 $layer=POLY_cond $X=4.27 $Y=1.557
+ $X2=4.305 $Y2=1.557
r51 20 21 59.2623 $w=3.66e-07 $l=4.5e-07 $layer=POLY_cond $X=3.82 $Y=1.557
+ $X2=4.27 $Y2=1.557
r52 19 20 1.97541 $w=3.66e-07 $l=1.5e-08 $layer=POLY_cond $X=3.805 $Y=1.557
+ $X2=3.82 $Y2=1.557
r53 16 25 3.88615 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.415 $Y2=1.565
r54 15 25 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.415 $Y2=1.565
r55 11 22 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.305 $Y=1.35
+ $X2=4.305 $Y2=1.557
r56 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.305 $Y=1.35
+ $X2=4.305 $Y2=0.74
r57 8 21 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.27 $Y=1.765
+ $X2=4.27 $Y2=1.557
r58 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.27 $Y=1.765
+ $X2=4.27 $Y2=2.4
r59 5 20 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.82 $Y=1.765
+ $X2=3.82 $Y2=1.557
r60 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.82 $Y=1.765
+ $X2=3.82 $Y2=2.4
r61 1 19 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.805 $Y=1.35
+ $X2=3.805 $Y2=1.557
r62 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.805 $Y=1.35
+ $X2=3.805 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%A_28_368# 1 2 3 10 12 14 16 19 20 21 24
c46 21 0 9.04372e-20 $X=1.4 $Y=2.99
r47 22 24 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=2.135 $Y=2.905
+ $X2=2.135 $Y2=2.375
r48 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.97 $Y=2.99
+ $X2=2.135 $Y2=2.905
r49 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.97 $Y=2.99 $X2=1.4
+ $Y2=2.99
r50 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.4 $Y2=2.99
r51 17 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.235 $Y2=2.815
r52 16 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.035
r53 16 19 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.815
r54 15 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.37 $Y=2.035
+ $X2=0.245 $Y2=2.035
r55 14 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=2.035
+ $X2=1.235 $Y2=2.035
r56 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.07 $Y=2.035 $X2=0.37
+ $Y2=2.035
r57 10 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.035
r58 10 12 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.815
r59 3 24 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.985
+ $Y=1.84 $X2=2.135 $Y2=2.375
r60 2 29 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.84 $X2=1.235 $Y2=2.115
r61 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.84 $X2=1.235 $Y2=2.815
r62 1 27 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r63 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
c50 13 0 1.88367e-19 $X=4.045 $Y=2.455
r51 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r53 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r54 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 27 30 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=0.735 $Y2=3.33
r59 25 27 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.735 $Y2=3.33
r63 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 18 31 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r65 18 28 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 16 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.88 $Y=3.33 $X2=3.6
+ $Y2=3.33
r67 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=4.005 $Y2=3.33
r68 15 33 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.13 $Y=3.33
+ $X2=4.56 $Y2=3.33
r69 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.13 $Y=3.33
+ $X2=4.005 $Y2=3.33
r70 11 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.005 $Y=3.245
+ $X2=4.005 $Y2=3.33
r71 11 13 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.005 $Y=3.245
+ $X2=4.005 $Y2=2.455
r72 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r73 7 9 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.455
r74 2 13 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.895
+ $Y=1.84 $X2=4.045 $Y2=2.455
r75 1 9 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%Y 1 2 3 4 15 17 18 23 25 27 31 34 37 40 43
r72 40 41 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=1.885
+ $X2=2.16 $Y2=2.035
r73 39 43 25.3036 $w=2.28e-07 $l=5.05e-07 $layer=LI1_cond $X=2.16 $Y=1.8
+ $X2=2.16 $Y2=1.295
r74 39 40 4.25903 $w=2.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.8 $X2=2.16
+ $Y2=1.885
r75 37 43 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.18
+ $X2=2.16 $Y2=1.295
r76 29 31 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=3.185 $Y=1.97
+ $X2=3.185 $Y2=1.985
r77 28 40 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.275 $Y=1.885
+ $X2=2.16 $Y2=1.885
r78 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.06 $Y=1.885
+ $X2=3.185 $Y2=1.97
r79 27 28 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.06 $Y=1.885
+ $X2=2.275 $Y2=1.885
r80 26 34 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.8 $Y=2.035
+ $X2=1.685 $Y2=2.035
r81 25 41 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.16 $Y2=2.035
r82 25 26 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=1.8 $Y2=2.035
r83 21 37 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=1.095
+ $X2=2.16 $Y2=1.095
r84 21 23 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.78 $Y=1.01
+ $X2=1.78 $Y2=0.76
r85 17 21 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=1.095
+ $X2=1.78 $Y2=1.095
r86 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.095
+ $X2=0.945 $Y2=1.095
r87 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.945 $Y2=1.095
r88 13 15 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.78 $Y2=0.76
r89 4 31 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.995
+ $Y=1.84 $X2=3.145 $Y2=1.985
r90 3 34 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=1.84 $X2=1.685 $Y2=2.115
r91 2 23 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.76
r92 1 15 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%A_510_368# 1 2 3 12 14 15 16 19 20 22 24
r45 22 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=2.12
+ $X2=4.495 $Y2=2.035
r46 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.495 $Y=2.12
+ $X2=4.495 $Y2=2.815
r47 21 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=2.035
+ $X2=3.595 $Y2=2.035
r48 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=2.035
+ $X2=4.495 $Y2=2.035
r49 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.33 $Y=2.035
+ $X2=3.68 $Y2=2.035
r50 17 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.595 $Y=2.905
+ $X2=3.595 $Y2=2.815
r51 16 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=2.12
+ $X2=3.595 $Y2=2.035
r52 16 19 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.595 $Y=2.12
+ $X2=3.595 $Y2=2.815
r53 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.51 $Y=2.99
+ $X2=3.595 $Y2=2.905
r54 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.51 $Y=2.99
+ $X2=2.86 $Y2=2.99
r55 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.695 $Y=2.905
+ $X2=2.86 $Y2=2.99
r56 10 12 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=2.695 $Y=2.905
+ $X2=2.695 $Y2=2.305
r57 3 29 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.84 $X2=4.495 $Y2=2.115
r58 3 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.84 $X2=4.495 $Y2=2.815
r59 2 27 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.595 $Y2=2.115
r60 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.595 $Y2=2.815
r61 1 12 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=2.55
+ $Y=1.84 $X2=2.695 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%A_27_74# 1 2 3 4 5 18 20 21 24 26 28 32 34
+ 38 40 45 47
r78 43 45 9.85637 $w=5.57e-07 $l=5.57225e-07 $layer=LI1_cond $X=2.45 $Y=0.515
+ $X2=2.69 $Y2=0.965
r79 41 43 3.83303 $w=5.57e-07 $l=1.75e-07 $layer=LI1_cond $X=2.45 $Y=0.34
+ $X2=2.45 $Y2=0.515
r80 36 38 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=4.56 $Y=1.01
+ $X2=4.56 $Y2=0.515
r81 35 47 7.02821 $w=1.7e-07 $l=1.36931e-07 $layer=LI1_cond $X=3.755 $Y=1.095
+ $X2=3.63 $Y2=1.07
r82 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.435 $Y=1.095
+ $X2=4.56 $Y2=1.01
r83 34 35 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.435 $Y=1.095
+ $X2=3.755 $Y2=1.095
r84 30 47 0.00168595 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=3.63 $Y=0.96
+ $X2=3.63 $Y2=1.07
r85 30 32 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.63 $Y=0.96
+ $X2=3.63 $Y2=0.515
r86 29 45 1.75224 $w=5.57e-07 $l=1.28938e-07 $layer=LI1_cond $X=2.785 $Y=1.045
+ $X2=2.69 $Y2=0.965
r87 28 47 7.02821 $w=1.7e-07 $l=1.36931e-07 $layer=LI1_cond $X=3.505 $Y=1.045
+ $X2=3.63 $Y2=1.07
r88 28 29 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.505 $Y=1.045
+ $X2=2.785 $Y2=1.045
r89 27 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0.34
+ $X2=1.28 $Y2=0.34
r90 26 41 7.83987 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.115 $Y=0.34
+ $X2=2.45 $Y2=0.34
r91 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=0.34
+ $X2=1.445 $Y2=0.34
r92 22 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.425
+ $X2=1.28 $Y2=0.34
r93 22 24 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.28 $Y=0.425
+ $X2=1.28 $Y2=0.675
r94 20 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0.34
+ $X2=1.28 $Y2=0.34
r95 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=0.34
+ $X2=0.445 $Y2=0.34
r96 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.445 $Y2=0.34
r97 16 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=0.425 $X2=0.28
+ $Y2=0.515
r98 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.38
+ $Y=0.37 $X2=4.52 $Y2=0.515
r99 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.45
+ $Y=0.37 $X2=3.59 $Y2=0.515
r100 3 45 121.333 $w=1.7e-07 $l=8.67929e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.69 $Y2=0.965
r101 3 43 121.333 $w=1.7e-07 $l=6.88694e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.69 $Y2=0.515
r102 2 24 182 $w=1.7e-07 $l=3.8461e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.37 $X2=1.28 $Y2=0.675
r103 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_2%VGND 1 2 9 13 15 17 25 32 33 36 39
r50 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r53 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r54 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=4.09
+ $Y2=0
r55 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=4.56
+ $Y2=0
r56 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r57 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r58 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r59 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=0 $X2=3.12
+ $Y2=0
r60 26 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.285 $Y=0 $X2=3.6
+ $Y2=0
r61 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=4.09
+ $Y2=0
r62 25 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.6
+ $Y2=0
r63 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r64 23 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r65 19 23 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r66 19 20 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r67 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=3.12
+ $Y2=0
r68 17 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=2.64
+ $Y2=0
r69 15 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r70 15 20 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=0.24
+ $Y2=0
r71 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0
r72 11 13 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0.675
r73 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=0.085 $X2=3.12
+ $Y2=0
r74 7 9 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.12 $Y=0.085 $X2=3.12
+ $Y2=0.625
r75 2 13 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=3.88
+ $Y=0.37 $X2=4.09 $Y2=0.675
r76 1 9 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.98
+ $Y=0.37 $X2=3.12 $Y2=0.625
.ends

