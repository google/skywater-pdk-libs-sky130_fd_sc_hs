# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__and3b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__and3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.260000 0.550000 1.930000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.440000 2.450000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.690000 1.350000 3.235000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.560000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.350000 3.715000 1.130000 ;
        RECT 3.410000 1.130000 3.715000 1.820000 ;
        RECT 3.410000 1.820000 3.755000 2.070000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.420000 0.375000 0.920000 ;
      RECT 0.115000  0.920000 1.230000 1.090000 ;
      RECT 0.115000  2.100000 1.070000 2.270000 ;
      RECT 0.115000  2.270000 0.400000 2.980000 ;
      RECT 0.545000  0.085000 0.875000 0.750000 ;
      RECT 0.570000  2.440000 0.900000 3.245000 ;
      RECT 0.900000  1.090000 1.230000 1.855000 ;
      RECT 0.900000  1.855000 1.070000 2.100000 ;
      RECT 1.400000  0.350000 1.755000 1.950000 ;
      RECT 1.400000  1.950000 2.750000 2.120000 ;
      RECT 1.400000  2.120000 1.730000 2.860000 ;
      RECT 1.900000  2.290000 2.230000 3.245000 ;
      RECT 2.420000  2.120000 2.750000 2.240000 ;
      RECT 2.420000  2.240000 4.215000 2.410000 ;
      RECT 2.420000  2.410000 2.750000 2.860000 ;
      RECT 2.815000  0.085000 3.145000 1.130000 ;
      RECT 2.960000  2.580000 3.290000 3.245000 ;
      RECT 3.875000  2.580000 4.205000 3.245000 ;
      RECT 3.885000  1.300000 4.215000 1.630000 ;
      RECT 3.895000  0.085000 4.145000 1.130000 ;
      RECT 4.045000  1.630000 4.215000 2.240000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__and3b_2
