* File: sky130_fd_sc_hs__or4bb_4.pex.spice
* Created: Thu Aug 27 21:07:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__OR4BB_4%D_N 3 5 7 8 12
c35 12 0 1.27147e-19 $X=0.59 $Y=1.515
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.515 $X2=0.59 $Y2=1.515
r37 8 12 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.515
r38 5 11 51.8789 $w=3.07e-07 $l=2.87228e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.585 $Y2=1.515
r39 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.34
r40 1 11 38.5336 $w=3.07e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.585 $Y2=1.515
r41 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%A_193_277# 1 2 3 10 12 13 15 16 18 19 21 22
+ 23 24 26 27 29 30 32 34 35 37 42 51 52 53 57 58 59 67 68 72 75 78
c181 35 0 7.31658e-20 $X=2.895 $Y=1.235
c182 32 0 1.39056e-19 $X=2.78 $Y=1.765
c183 27 0 1.38753e-19 $X=2.09 $Y=1.235
c184 13 0 2.40437e-20 $X=1.07 $Y=1.235
c185 10 0 1.27147e-19 $X=1.055 $Y=1.765
r186 77 78 12.3324 $w=9.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=0.805
+ $X2=6.28 $Y2=0.805
r187 74 77 0.737363 $w=9.08e-07 $l=5.5e-08 $layer=LI1_cond $X=6.06 $Y=0.805
+ $X2=6.115 $Y2=0.805
r188 74 75 1.60122 $w=9.08e-07 $l=8.5e-08 $layer=LI1_cond $X=6.06 $Y=0.805
+ $X2=5.975 $Y2=0.805
r189 70 72 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=7.19 $Y=1.09
+ $X2=7.19 $Y2=0.515
r190 68 70 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.025 $Y=1.175
+ $X2=7.19 $Y2=1.09
r191 68 78 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.025 $Y=1.175
+ $X2=6.28 $Y2=1.175
r192 66 74 11.0791 $w=1.7e-07 $l=4.55e-07 $layer=LI1_cond $X=6.06 $Y=1.26
+ $X2=6.06 $Y2=0.805
r193 66 67 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.06 $Y=1.26 $X2=6.06
+ $Y2=1.76
r194 65 75 3.95999 $w=7.38e-07 $l=2.45e-07 $layer=LI1_cond $X=5.73 $Y=0.72
+ $X2=5.975 $Y2=0.72
r195 62 65 12.6073 $w=7.38e-07 $l=7.8e-07 $layer=LI1_cond $X=4.95 $Y=0.72
+ $X2=5.73 $Y2=0.72
r196 58 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.975 $Y=1.845
+ $X2=6.06 $Y2=1.76
r197 58 59 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=5.975 $Y=1.845
+ $X2=4.715 $Y2=1.845
r198 55 57 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.55 $Y=2.29 $X2=4.55
+ $Y2=2.2
r199 54 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.55 $Y=1.93
+ $X2=4.715 $Y2=1.845
r200 54 57 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.55 $Y=1.93
+ $X2=4.55 $Y2=2.2
r201 52 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.385 $Y=2.375
+ $X2=4.55 $Y2=2.29
r202 52 53 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=4.385 $Y=2.375
+ $X2=3.205 $Y2=2.375
r203 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.12 $Y=2.29
+ $X2=3.205 $Y2=2.375
r204 50 51 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.12 $Y=1.54
+ $X2=3.12 $Y2=2.29
r205 44 48 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.125 $Y=1.4
+ $X2=2.805 $Y2=1.4
r206 42 50 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.035 $Y=1.4
+ $X2=3.12 $Y2=1.54
r207 42 48 9.4665 $w=2.78e-07 $l=2.3e-07 $layer=LI1_cond $X=3.035 $Y=1.4
+ $X2=2.805 $Y2=1.4
r208 40 41 0.551487 $w=4.37e-07 $l=5e-09 $layer=POLY_cond $X=1.5 $Y=1.5
+ $X2=1.505 $Y2=1.5
r209 39 40 47.4279 $w=4.37e-07 $l=4.3e-07 $layer=POLY_cond $X=1.07 $Y=1.5
+ $X2=1.5 $Y2=1.5
r210 38 39 1.65446 $w=4.37e-07 $l=1.5e-08 $layer=POLY_cond $X=1.055 $Y=1.5
+ $X2=1.07 $Y2=1.5
r211 35 37 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.895 $Y=1.235
+ $X2=2.895 $Y2=0.74
r212 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.78 $Y=1.765
+ $X2=2.78 $Y2=2.4
r213 30 32 79.6222 $w=2.42e-07 $l=3.89198e-07 $layer=POLY_cond $X=2.83 $Y=1.4
+ $X2=2.78 $Y2=1.765
r214 30 35 39.7875 $w=2.42e-07 $l=1.94808e-07 $layer=POLY_cond $X=2.83 $Y=1.4
+ $X2=2.895 $Y2=1.235
r215 30 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.4 $X2=2.805 $Y2=1.4
r216 27 29 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.09 $Y=1.235
+ $X2=2.09 $Y2=0.74
r217 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.05 $Y=1.765
+ $X2=2.05 $Y2=2.4
r218 23 41 12.929 $w=4.37e-07 $l=1.3784e-07 $layer=POLY_cond $X=1.595 $Y=1.4
+ $X2=1.505 $Y2=1.5
r219 22 24 92.9106 $w=1.95e-07 $l=3.70951e-07 $layer=POLY_cond $X=2.062 $Y=1.4
+ $X2=2.05 $Y2=1.765
r220 22 27 43.4747 $w=1.95e-07 $l=1.78452e-07 $layer=POLY_cond $X=2.062 $Y=1.4
+ $X2=2.09 $Y2=1.235
r221 22 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.4 $X2=2.125 $Y2=1.4
r222 22 30 91.8022 $w=3.3e-07 $l=5.25e-07 $layer=POLY_cond $X=2.165 $Y=1.4
+ $X2=2.69 $Y2=1.4
r223 22 23 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=1.96 $Y=1.4
+ $X2=1.595 $Y2=1.4
r224 19 41 28.039 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.5
r225 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r226 16 40 28.039 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.5 $Y=1.235
+ $X2=1.5 $Y2=1.5
r227 16 18 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.5 $Y=1.235
+ $X2=1.5 $Y2=0.74
r228 13 39 28.039 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.07 $Y=1.235
+ $X2=1.07 $Y2=1.5
r229 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.07 $Y=1.235
+ $X2=1.07 $Y2=0.74
r230 10 38 28.039 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=1.5
r231 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=2.4
r232 3 57 600 $w=1.7e-07 $l=3.05941e-07 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.96 $X2=4.55 $Y2=2.2
r233 2 72 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.05
+ $Y=0.37 $X2=7.19 $Y2=0.515
r234 1 77 91 $w=1.7e-07 $l=1.37559e-06 $layer=licon1_NDIFF $count=2 $X=4.81
+ $Y=0.37 $X2=6.115 $Y2=0.515
r235 1 65 60.6667 $w=1.7e-07 $l=9.89848e-07 $layer=licon1_NDIFF $count=3 $X=4.81
+ $Y=0.37 $X2=5.73 $Y2=0.515
r236 1 62 60.6667 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=3 $X=4.81
+ $Y=0.37 $X2=4.95 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%C_N 1 3 6 8 12
c37 12 0 1.39056e-19 $X=3.54 $Y=1.515
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.54
+ $Y=1.515 $X2=3.54 $Y2=1.515
r39 8 12 5.08431 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=3.545 $Y=1.665
+ $X2=3.545 $Y2=1.515
r40 4 11 39.9551 $w=4.18e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.405 $Y=1.35
+ $X2=3.465 $Y2=1.515
r41 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.405 $Y=1.35
+ $X2=3.405 $Y2=0.79
r42 1 11 49.7565 $w=4.18e-07 $l=3.16228e-07 $layer=POLY_cond $X=3.315 $Y=1.765
+ $X2=3.465 $Y2=1.515
r43 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.765
+ $X2=3.315 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%A_27_94# 1 2 8 9 11 12 14 16 17 19 22 27 28
+ 29 31 32 33 34 35 37 38 40 41 42
r145 46 49 27.2711 $w=3.8e-07 $l=2.15e-07 $layer=POLY_cond $X=4.11 $Y=1.195
+ $X2=4.325 $Y2=1.195
r146 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.11
+ $Y=1.085 $X2=4.11 $Y2=1.085
r147 42 45 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.11 $Y=1.005 $X2=4.11
+ $Y2=1.085
r148 40 41 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.115
+ $X2=0.265 $Y2=1.95
r149 38 41 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.17 $Y=1.13
+ $X2=0.17 $Y2=1.95
r150 36 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.78 $Y=1.88
+ $X2=2.78 $Y2=2.39
r151 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.695 $Y=1.795
+ $X2=2.78 $Y2=1.88
r152 34 35 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.695 $Y=1.795
+ $X2=1.79 $Y2=1.795
r153 32 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=1.005
+ $X2=4.11 $Y2=1.005
r154 32 33 140.594 $w=1.68e-07 $l=2.155e-06 $layer=LI1_cond $X=3.945 $Y=1.005
+ $X2=1.79 $Y2=1.005
r155 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=1.71
+ $X2=1.79 $Y2=1.795
r156 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=1.09
+ $X2=1.79 $Y2=1.005
r157 30 31 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.705 $Y=1.09
+ $X2=1.705 $Y2=1.71
r158 28 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.695 $Y=2.475
+ $X2=2.78 $Y2=2.39
r159 28 29 146.791 $w=1.68e-07 $l=2.25e-06 $layer=LI1_cond $X=2.695 $Y=2.475
+ $X2=0.445 $Y2=2.475
r160 27 29 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.265 $Y=2.39
+ $X2=0.445 $Y2=2.475
r161 26 40 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.115
r162 26 27 8.3232 $w=3.58e-07 $l=2.6e-07 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.39
r163 20 38 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=1.13
r164 20 22 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.615
r165 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.885
+ $X2=4.775 $Y2=2.46
r166 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.775 $Y=1.795
+ $X2=4.775 $Y2=1.885
r167 15 51 20.2441 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=4.775 $Y=1.47
+ $X2=4.775 $Y2=1.195
r168 15 16 126.331 $w=1.8e-07 $l=3.25e-07 $layer=POLY_cond $X=4.775 $Y=1.47
+ $X2=4.775 $Y2=1.795
r169 12 51 5.07368 $w=3.8e-07 $l=4e-08 $layer=POLY_cond $X=4.735 $Y=1.195
+ $X2=4.775 $Y2=1.195
r170 12 49 52.0053 $w=3.8e-07 $l=4.1e-07 $layer=POLY_cond $X=4.735 $Y=1.195
+ $X2=4.325 $Y2=1.195
r171 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.735 $Y=1.185
+ $X2=4.735 $Y2=0.74
r172 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.325 $Y=1.885
+ $X2=4.325 $Y2=2.46
r173 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.325 $Y=1.795
+ $X2=4.325 $Y2=1.885
r174 7 49 20.2441 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=4.325 $Y=1.47
+ $X2=4.325 $Y2=1.195
r175 7 8 126.331 $w=1.8e-07 $l=3.25e-07 $layer=POLY_cond $X=4.325 $Y=1.47
+ $X2=4.325 $Y2=1.795
r176 2 40 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r177 1 22 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.47 $X2=0.28 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%A_678_368# 1 2 8 9 11 13 14 16 17 21 23 27
+ 30 31 32 34 37 43 44 49
c101 43 0 7.31658e-20 $X=3.785 $Y=0.6
r102 48 49 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.725 $Y=1.425
+ $X2=5.815 $Y2=1.425
r103 41 43 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0.6
+ $X2=3.785 $Y2=0.6
r104 38 48 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.64 $Y=1.425
+ $X2=5.725 $Y2=1.425
r105 38 45 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=5.64 $Y=1.425
+ $X2=5.225 $Y2=1.425
r106 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.64
+ $Y=1.425 $X2=5.64 $Y2=1.425
r107 35 44 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.615 $Y=1.425
+ $X2=4.53 $Y2=1.425
r108 35 37 35.7956 $w=3.28e-07 $l=1.025e-06 $layer=LI1_cond $X=4.615 $Y=1.425
+ $X2=5.64 $Y2=1.425
r109 34 44 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.53 $Y=1.26
+ $X2=4.53 $Y2=1.425
r110 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.53 $Y=0.75
+ $X2=4.53 $Y2=1.26
r111 31 44 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.445 $Y=1.505
+ $X2=4.53 $Y2=1.425
r112 31 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.445 $Y=1.505
+ $X2=4.055 $Y2=1.505
r113 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.97 $Y=1.59
+ $X2=4.055 $Y2=1.505
r114 29 30 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.97 $Y=1.59
+ $X2=3.97 $Y2=1.95
r115 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.445 $Y=0.665
+ $X2=4.53 $Y2=0.75
r116 27 43 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.445 $Y=0.665
+ $X2=3.785 $Y2=0.665
r117 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.885 $Y=2.035
+ $X2=3.97 $Y2=1.95
r118 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.885 $Y=2.035
+ $X2=3.54 $Y2=2.035
r119 19 21 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.33 $Y=1.26
+ $X2=6.33 $Y2=0.74
r120 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.255 $Y=1.335
+ $X2=6.33 $Y2=1.26
r121 17 49 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.255 $Y=1.335
+ $X2=5.815 $Y2=1.335
r122 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.725 $Y=1.885
+ $X2=5.725 $Y2=2.46
r123 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.725 $Y=1.795
+ $X2=5.725 $Y2=1.885
r124 12 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=1.59
+ $X2=5.725 $Y2=1.425
r125 12 13 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=5.725 $Y=1.59
+ $X2=5.725 $Y2=1.795
r126 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.225 $Y=1.885
+ $X2=5.225 $Y2=2.46
r127 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.225 $Y=1.795
+ $X2=5.225 $Y2=1.885
r128 7 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.225 $Y=1.59
+ $X2=5.225 $Y2=1.425
r129 7 8 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=5.225 $Y=1.59
+ $X2=5.225 $Y2=1.795
r130 2 25 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.84 $X2=3.54 $Y2=2.035
r131 1 41 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=3.48
+ $Y=0.47 $X2=3.62 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%B 1 3 6 8 10 11 12 19
c55 1 0 8.95903e-20 $X=6.735 $Y=1.885
r56 19 20 25.9538 $w=3.9e-07 $l=2.1e-07 $layer=POLY_cond $X=6.975 $Y=1.667
+ $X2=7.185 $Y2=1.667
r57 17 19 20.3923 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=6.81 $Y=1.667
+ $X2=6.975 $Y2=1.667
r58 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.81
+ $Y=1.615 $X2=6.81 $Y2=1.615
r59 15 17 9.26923 $w=3.9e-07 $l=7.5e-08 $layer=POLY_cond $X=6.735 $Y=1.667
+ $X2=6.81 $Y2=1.667
r60 12 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.96 $Y=1.615
+ $X2=6.81 $Y2=1.615
r61 11 18 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.81 $Y2=1.615
r62 8 20 25.2441 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.185 $Y=1.885
+ $X2=7.185 $Y2=1.667
r63 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.185 $Y=1.885
+ $X2=7.185 $Y2=2.46
r64 4 19 25.2441 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.975 $Y=1.45
+ $X2=6.975 $Y2=1.667
r65 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.975 $Y=1.45
+ $X2=6.975 $Y2=0.74
r66 1 15 25.2441 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.735 $Y=1.885
+ $X2=6.735 $Y2=1.667
r67 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.735 $Y=1.885
+ $X2=6.735 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%A 1 3 5 6 8 10 11 13 14 15 26
c46 11 0 9.04372e-20 $X=8.135 $Y=1.885
c47 6 0 4.65189e-20 $X=7.635 $Y=1.885
r48 26 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.37
+ $Y=1.385 $X2=8.37 $Y2=1.385
r49 24 26 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=8.135 $Y=1.385
+ $X2=8.37 $Y2=1.385
r50 22 24 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=7.69 $Y=1.385
+ $X2=8.135 $Y2=1.385
r51 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.69
+ $Y=1.385 $X2=7.69 $Y2=1.385
r52 20 22 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=7.635 $Y=1.385
+ $X2=7.69 $Y2=1.385
r53 18 20 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=7.59 $Y=1.385
+ $X2=7.635 $Y2=1.385
r54 15 27 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=8.4 $Y=1.365 $X2=8.37
+ $Y2=1.365
r55 14 27 14.0162 $w=3.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.92 $Y=1.365
+ $X2=8.37 $Y2=1.365
r56 14 23 7.16384 $w=3.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.92 $Y=1.365
+ $X2=7.69 $Y2=1.365
r57 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.135 $Y=1.885
+ $X2=8.135 $Y2=2.46
r58 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.135 $Y=1.795
+ $X2=8.135 $Y2=1.885
r59 9 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.135 $Y=1.55
+ $X2=8.135 $Y2=1.385
r60 9 10 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=8.135 $Y=1.55
+ $X2=8.135 $Y2=1.795
r61 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.635 $Y=1.885
+ $X2=7.635 $Y2=2.46
r62 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.635 $Y=1.795 $X2=7.635
+ $Y2=1.885
r63 4 20 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.635 $Y=1.55
+ $X2=7.635 $Y2=1.385
r64 4 5 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=7.635 $Y=1.55
+ $X2=7.635 $Y2=1.795
r65 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.59 $Y=1.22
+ $X2=7.59 $Y2=1.385
r66 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.59 $Y=1.22 $X2=7.59
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%VPWR 1 2 3 4 17 21 25 29 31 33 38 43 50 51
+ 54 57 60 63
r83 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r84 60 61 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r86 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 51 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r88 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r89 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=3.33
+ $X2=7.91 $Y2=3.33
r90 48 50 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=3.33
+ $X2=8.4 $Y2=3.33
r91 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r92 46 47 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r93 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=3.33
+ $X2=3.005 $Y2=3.33
r94 44 46 278.578 $w=1.68e-07 $l=4.27e-06 $layer=LI1_cond $X=3.17 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=3.33
+ $X2=7.91 $Y2=3.33
r96 43 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=3.33
+ $X2=7.44 $Y2=3.33
r97 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r98 42 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 39 57 10.2049 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=1.99 $Y=3.33
+ $X2=1.777 $Y2=3.33
r101 39 41 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.99 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=3.33
+ $X2=3.005 $Y2=3.33
r103 38 41 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.84 $Y=3.33 $X2=2.64
+ $Y2=3.33
r104 37 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r105 37 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r106 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r107 34 54 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.822 $Y2=3.33
r108 34 36 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 33 57 10.2049 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.777 $Y2=3.33
r110 33 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 31 47 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 31 61 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 27 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=3.245
+ $X2=7.91 $Y2=3.33
r114 27 29 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=7.91 $Y=3.245
+ $X2=7.91 $Y2=2.495
r115 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=3.245
+ $X2=3.005 $Y2=3.33
r116 23 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.005 $Y=3.245
+ $X2=3.005 $Y2=2.815
r117 19 57 1.63918 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.777 $Y=3.245
+ $X2=1.777 $Y2=3.33
r118 19 21 11.66 $w=4.23e-07 $l=4.3e-07 $layer=LI1_cond $X=1.777 $Y=3.245
+ $X2=1.777 $Y2=2.815
r119 15 54 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.822 $Y=3.245
+ $X2=0.822 $Y2=3.33
r120 15 17 14.3638 $w=3.43e-07 $l=4.3e-07 $layer=LI1_cond $X=0.822 $Y=3.245
+ $X2=0.822 $Y2=2.815
r121 4 29 300 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=2 $X=7.71
+ $Y=1.96 $X2=7.91 $Y2=2.495
r122 3 25 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.84 $X2=3.005 $Y2=2.815
r123 2 21 600 $w=1.7e-07 $l=1.06806e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.775 $Y2=2.815
r124 1 17 600 $w=1.7e-07 $l=1.0884e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.82 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%X 1 2 3 4 19 21 26 29 30 31 32 39 47 49
c54 47 0 1.38753e-19 $X=1.267 $Y=1.18
c55 29 0 2.40437e-20 $X=2.14 $Y=0.585
r56 38 49 2.11544 $w=3.63e-07 $l=6.7e-08 $layer=LI1_cond $X=1.267 $Y=1.362
+ $X2=1.267 $Y2=1.295
r57 32 39 2.55837 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.267 $Y=2.135
+ $X2=1.267 $Y2=2.05
r58 32 39 1.57869 $w=3.63e-07 $l=5e-08 $layer=LI1_cond $X=1.267 $Y=2 $X2=1.267
+ $Y2=2.05
r59 31 32 10.5772 $w=3.63e-07 $l=3.35e-07 $layer=LI1_cond $X=1.267 $Y=1.665
+ $X2=1.267 $Y2=2
r60 30 49 0.284164 $w=3.63e-07 $l=9e-09 $layer=LI1_cond $X=1.267 $Y=1.286
+ $X2=1.267 $Y2=1.295
r61 30 47 3.47695 $w=3.63e-07 $l=1.06e-07 $layer=LI1_cond $X=1.267 $Y=1.286
+ $X2=1.267 $Y2=1.18
r62 30 31 9.28269 $w=3.63e-07 $l=2.94e-07 $layer=LI1_cond $X=1.267 $Y=1.371
+ $X2=1.267 $Y2=1.665
r63 30 38 0.284164 $w=3.63e-07 $l=9e-09 $layer=LI1_cond $X=1.267 $Y=1.371
+ $X2=1.267 $Y2=1.362
r64 26 28 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.285 $Y=0.515
+ $X2=1.285 $Y2=0.665
r65 21 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.585
+ $X2=2.14 $Y2=0.585
r66 21 23 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.305 $Y=0.585
+ $X2=2.68 $Y2=0.585
r67 17 32 5.50802 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=1.45 $Y=2.135
+ $X2=1.267 $Y2=2.135
r68 17 19 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.45 $Y=2.135
+ $X2=2.315 $Y2=2.135
r69 16 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0.665
+ $X2=1.285 $Y2=0.665
r70 16 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.45 $Y=0.665
+ $X2=2.14 $Y2=0.665
r71 13 28 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.75
+ $X2=1.285 $Y2=0.665
r72 13 47 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.285 $Y=0.75
+ $X2=1.285 $Y2=1.18
r73 4 19 600 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=1.84 $X2=2.315 $Y2=2.135
r74 3 32 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.84 $X2=1.28 $Y2=2.02
r75 2 23 91 $w=1.7e-07 $l=6.13148e-07 $layer=licon1_NDIFF $count=2 $X=2.165
+ $Y=0.37 $X2=2.68 $Y2=0.585
r76 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.145
+ $Y=0.37 $X2=1.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%A_791_392# 1 2 3 14 18 22 23
r34 21 23 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=2.852
+ $X2=5.165 $Y2=2.852
r35 21 22 4.83021 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=2.852
+ $X2=4.835 $Y2=2.852
r36 16 18 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=5.99 $Y=2.905 $X2=5.99
+ $Y2=2.605
r37 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.865 $Y=2.99
+ $X2=5.99 $Y2=2.905
r38 14 23 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.865 $Y=2.99
+ $X2=5.165 $Y2=2.99
r39 12 22 24.2013 $w=3.48e-07 $l=7.35e-07 $layer=LI1_cond $X=4.1 $Y=2.805
+ $X2=4.835 $Y2=2.805
r40 3 18 600 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.96 $X2=5.95 $Y2=2.605
r41 2 21 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=4.85
+ $Y=1.96 $X2=5 $Y2=2.805
r42 1 12 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=3.955
+ $Y=1.96 $X2=4.1 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%A_1060_392# 1 2 13 16 18 19
r30 18 19 16.3833 $w=3.18e-07 $l=3.85e-07 $layer=LI1_cond $X=6.96 $Y=2.11
+ $X2=6.575 $Y2=2.11
r31 11 18 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.96 $Y=2.27 $X2=6.96
+ $Y2=2.11
r32 11 13 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.96 $Y=2.27 $X2=6.96
+ $Y2=2.57
r33 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=2.185
+ $X2=5.5 $Y2=2.185
r34 10 19 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=5.665 $Y=2.185
+ $X2=6.575 $Y2=2.185
r35 2 18 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.96 $X2=6.96 $Y2=2.115
r36 2 13 600 $w=1.7e-07 $l=6.80882e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.96 $X2=6.96 $Y2=2.57
r37 1 16 300 $w=1.7e-07 $l=3.09233e-07 $layer=licon1_PDIFF $count=2 $X=5.3
+ $Y=1.96 $X2=5.5 $Y2=2.185
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%A_1273_392# 1 2 3 12 14 15 16 19 20 22 24
c53 22 0 4.65189e-20 $X=8.387 $Y=2.24
c54 16 0 8.95903e-20 $X=7.41 $Y=2.24
c55 14 0 9.04372e-20 $X=7.245 $Y=2.99
r56 22 29 3.48019 $w=2.75e-07 $l=1.62942e-07 $layer=LI1_cond $X=8.387 $Y=2.24
+ $X2=8.36 $Y2=2.09
r57 22 24 9.01001 $w=2.73e-07 $l=2.15e-07 $layer=LI1_cond $X=8.387 $Y=2.24
+ $X2=8.387 $Y2=2.455
r58 21 27 3.64781 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.575 $Y=2.095
+ $X2=7.41 $Y2=2.095
r59 20 29 3.34255 $w=2.9e-07 $l=1.67481e-07 $layer=LI1_cond $X=8.195 $Y=2.095
+ $X2=8.36 $Y2=2.09
r60 20 21 24.6384 $w=2.88e-07 $l=6.2e-07 $layer=LI1_cond $X=8.195 $Y=2.095
+ $X2=7.575 $Y2=2.095
r61 17 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.41 $Y=2.905 $X2=7.41
+ $Y2=2.815
r62 16 27 3.20565 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=7.41 $Y=2.24
+ $X2=7.41 $Y2=2.095
r63 16 19 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=7.41 $Y=2.24
+ $X2=7.41 $Y2=2.815
r64 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.245 $Y=2.99
+ $X2=7.41 $Y2=2.905
r65 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.245 $Y=2.99
+ $X2=6.675 $Y2=2.99
r66 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.51 $Y=2.905
+ $X2=6.675 $Y2=2.99
r67 10 12 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=6.51 $Y=2.905 $X2=6.51
+ $Y2=2.605
r68 3 29 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.96 $X2=8.36 $Y2=2.105
r69 3 24 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=8.21
+ $Y=1.96 $X2=8.36 $Y2=2.455
r70 2 27 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.96 $X2=7.41 $Y2=2.115
r71 2 19 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.96 $X2=7.41 $Y2=2.815
r72 1 12 600 $w=1.7e-07 $l=7.13828e-07 $layer=licon1_PDIFF $count=1 $X=6.365
+ $Y=1.96 $X2=6.51 $Y2=2.605
.ends

.subckt PM_SKY130_FD_SC_HS__OR4BB_4%VGND 1 2 3 4 5 6 21 23 27 31 35 39 41 43 48
+ 53 60 61 64 68 74 79 85 87 90
r91 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r92 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r93 84 88 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r94 83 85 6.58698 $w=4.93e-07 $l=4.5e-08 $layer=LI1_cond $X=4.56 $Y=0.162
+ $X2=4.605 $Y2=0.162
r95 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r96 81 83 6.0408 $w=4.93e-07 $l=2.5e-07 $layer=LI1_cond $X=4.31 $Y=0.162
+ $X2=4.56 $Y2=0.162
r97 77 81 5.55754 $w=4.93e-07 $l=2.3e-07 $layer=LI1_cond $X=4.08 $Y=0.162
+ $X2=4.31 $Y2=0.162
r98 77 79 7.07024 $w=4.93e-07 $l=6.5e-08 $layer=LI1_cond $X=4.08 $Y=0.162
+ $X2=4.015 $Y2=0.162
r99 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r100 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r101 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r102 68 71 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=1.795 $Y2=0.325
r103 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r104 65 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r105 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r106 61 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r107 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r108 58 90 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.31 $Y=0 $X2=7.975
+ $Y2=0
r109 58 60 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.31 $Y=0 $X2=8.4
+ $Y2=0
r110 57 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r111 57 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r112 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r113 54 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=0 $X2=6.615
+ $Y2=0
r114 54 56 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.78 $Y=0 $X2=7.44
+ $Y2=0
r115 53 90 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.975
+ $Y2=0
r116 53 56 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.44
+ $Y2=0
r117 52 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r118 52 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r119 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r120 49 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.96 $Y=0 $X2=1.795
+ $Y2=0
r121 49 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.96 $Y=0 $X2=2.64
+ $Y2=0
r122 48 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.11
+ $Y2=0
r123 48 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.945 $Y=0
+ $X2=2.64 $Y2=0
r124 46 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r125 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r126 43 64 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.765
+ $Y2=0
r127 43 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r128 41 84 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r129 41 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r130 37 90 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.975 $Y=0.085
+ $X2=7.975 $Y2=0
r131 37 39 7.67632 $w=6.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.975 $Y=0.085
+ $X2=7.975 $Y2=0.515
r132 33 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.615 $Y=0.085
+ $X2=6.615 $Y2=0
r133 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.615 $Y=0.085
+ $X2=6.615 $Y2=0.495
r134 31 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.45 $Y=0 $X2=6.615
+ $Y2=0
r135 31 85 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=6.45 $Y=0
+ $X2=4.605 $Y2=0
r136 30 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.11
+ $Y2=0
r137 30 79 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.275 $Y=0
+ $X2=4.015 $Y2=0
r138 25 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=0.085
+ $X2=3.11 $Y2=0
r139 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.11 $Y=0.085
+ $X2=3.11 $Y2=0.55
r140 24 64 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.765
+ $Y2=0
r141 23 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.795
+ $Y2=0
r142 23 24 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.63 $Y=0
+ $X2=0.915 $Y2=0
r143 19 64 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0
r144 19 21 20.3598 $w=2.98e-07 $l=5.3e-07 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0.615
r145 6 39 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=7.665
+ $Y=0.37 $X2=8.145 $Y2=0.515
r146 5 35 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=6.405
+ $Y=0.37 $X2=6.615 $Y2=0.495
r147 4 81 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.18 $X2=4.31 $Y2=0.325
r148 3 27 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.97 $Y=0.37
+ $X2=3.11 $Y2=0.55
r149 2 71 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=1.575
+ $Y=0.37 $X2=1.795 $Y2=0.325
r150 1 21 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.47 $X2=0.78 $Y2=0.615
.ends

