# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__mux4_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__mux4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.215000 1.320000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.000000 1.215000 3.330000 2.150000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.500000 1.215000 3.870000 2.150000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.850000 1.445000 6.180000 1.780000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.738000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.450000 1.215000 0.820000 1.780000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.205000 1.350000 8.535000 1.780000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.558100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.080000 0.400000 9.485000 1.180000 ;
        RECT 9.220000 2.560000 9.485000 2.890000 ;
        RECT 9.245000 1.180000 9.485000 2.560000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
        RECT 0.700000  0.085000 1.090000 0.680000 ;
        RECT 3.125000  0.085000 3.715000 0.680000 ;
        RECT 5.260000  0.085000 5.590000 0.935000 ;
        RECT 8.580000  0.085000 8.910000 1.180000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.600000 3.415000 ;
        RECT 0.725000 1.950000 1.055000 3.245000 ;
        RECT 3.265000 2.675000 3.595000 3.245000 ;
        RECT 5.730000 2.675000 6.060000 3.245000 ;
        RECT 8.690000 2.290000 9.020000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.110000 0.350000 0.445000 0.860000 ;
      RECT 0.110000 0.860000 1.700000 1.030000 ;
      RECT 0.110000 1.030000 0.280000 1.950000 ;
      RECT 0.110000 1.950000 0.555000 2.880000 ;
      RECT 1.530000 0.255000 2.630000 0.425000 ;
      RECT 1.530000 0.425000 1.700000 0.860000 ;
      RECT 1.530000 1.030000 1.700000 1.200000 ;
      RECT 1.530000 1.200000 1.860000 1.530000 ;
      RECT 1.875000 0.595000 2.200000 1.030000 ;
      RECT 2.030000 1.030000 2.200000 1.685000 ;
      RECT 2.030000 1.685000 2.550000 2.335000 ;
      RECT 2.030000 2.335000 4.020000 2.505000 ;
      RECT 2.030000 2.505000 2.550000 2.725000 ;
      RECT 2.460000 0.425000 2.630000 0.875000 ;
      RECT 2.460000 0.875000 4.750000 1.045000 ;
      RECT 2.460000 1.045000 2.790000 1.450000 ;
      RECT 3.795000 2.505000 4.020000 2.905000 ;
      RECT 3.795000 2.905000 5.550000 3.075000 ;
      RECT 4.080000 1.045000 4.410000 1.450000 ;
      RECT 4.210000 0.375000 5.090000 0.705000 ;
      RECT 4.305000 1.995000 5.680000 2.165000 ;
      RECT 4.305000 2.165000 5.165000 2.735000 ;
      RECT 4.580000 1.045000 4.750000 1.445000 ;
      RECT 4.580000 1.445000 5.340000 1.775000 ;
      RECT 4.920000 0.705000 5.090000 1.105000 ;
      RECT 4.920000 1.105000 6.235000 1.275000 ;
      RECT 5.350000 2.335000 6.620000 2.505000 ;
      RECT 5.350000 2.505000 5.550000 2.905000 ;
      RECT 5.510000 1.275000 5.680000 1.995000 ;
      RECT 5.985000 0.265000 7.695000 0.435000 ;
      RECT 5.985000 0.435000 6.485000 0.445000 ;
      RECT 5.985000 0.445000 6.235000 1.105000 ;
      RECT 6.290000 1.950000 6.620000 2.335000 ;
      RECT 6.290000 2.505000 6.620000 2.980000 ;
      RECT 6.405000 0.615000 7.355000 0.785000 ;
      RECT 6.405000 0.785000 6.575000 1.950000 ;
      RECT 6.745000 0.955000 6.925000 1.115000 ;
      RECT 6.745000 1.115000 7.120000 1.285000 ;
      RECT 6.790000 1.285000 7.120000 2.905000 ;
      RECT 6.790000 2.905000 8.520000 3.075000 ;
      RECT 7.105000 0.605000 7.355000 0.615000 ;
      RECT 7.105000 0.785000 7.355000 0.935000 ;
      RECT 7.290000 1.105000 7.695000 1.275000 ;
      RECT 7.290000 1.275000 7.460000 1.945000 ;
      RECT 7.290000 1.945000 7.620000 2.735000 ;
      RECT 7.525000 0.435000 7.695000 1.105000 ;
      RECT 7.630000 1.445000 8.035000 1.775000 ;
      RECT 7.850000 1.775000 8.035000 1.950000 ;
      RECT 7.850000 1.950000 8.180000 2.735000 ;
      RECT 7.865000 0.500000 8.410000 1.180000 ;
      RECT 7.865000 1.180000 8.035000 1.445000 ;
      RECT 8.350000 1.950000 8.915000 2.120000 ;
      RECT 8.350000 2.120000 8.520000 2.905000 ;
      RECT 8.745000 1.350000 9.075000 1.680000 ;
      RECT 8.745000 1.680000 8.915000 1.950000 ;
  END
END sky130_fd_sc_hs__mux4_1
