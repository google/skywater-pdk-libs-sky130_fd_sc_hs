* File: sky130_fd_sc_hs__nand2b_4.pxi.spice
* Created: Thu Aug 27 20:50:47 2020
* 
x_PM_SKY130_FD_SC_HS__NAND2B_4%A_N N_A_N_M1012_g N_A_N_c_91_n N_A_N_M1005_g
+ N_A_N_c_86_n N_A_N_c_93_n N_A_N_M1008_g N_A_N_c_87_n N_A_N_c_88_n A_N A_N
+ N_A_N_c_89_n N_A_N_c_90_n PM_SKY130_FD_SC_HS__NAND2B_4%A_N
x_PM_SKY130_FD_SC_HS__NAND2B_4%A_31_74# N_A_31_74#_M1012_s N_A_31_74#_M1005_d
+ N_A_31_74#_c_138_n N_A_31_74#_M1000_g N_A_31_74#_c_139_n N_A_31_74#_c_140_n
+ N_A_31_74#_c_141_n N_A_31_74#_M1007_g N_A_31_74#_c_151_n N_A_31_74#_M1003_g
+ N_A_31_74#_c_142_n N_A_31_74#_M1010_g N_A_31_74#_c_152_n N_A_31_74#_M1006_g
+ N_A_31_74#_c_143_n N_A_31_74#_M1014_g N_A_31_74#_c_144_n N_A_31_74#_c_145_n
+ N_A_31_74#_c_146_n N_A_31_74#_c_153_n N_A_31_74#_c_147_n N_A_31_74#_c_148_n
+ N_A_31_74#_c_155_n N_A_31_74#_c_149_n N_A_31_74#_c_150_n
+ PM_SKY130_FD_SC_HS__NAND2B_4%A_31_74#
x_PM_SKY130_FD_SC_HS__NAND2B_4%B N_B_M1001_g N_B_c_256_n N_B_c_257_n N_B_M1004_g
+ N_B_M1009_g N_B_c_264_n N_B_M1002_g N_B_c_265_n N_B_M1013_g N_B_M1011_g B B B
+ N_B_c_262_n N_B_c_263_n N_B_c_288_p PM_SKY130_FD_SC_HS__NAND2B_4%B
x_PM_SKY130_FD_SC_HS__NAND2B_4%VPWR N_VPWR_M1005_s N_VPWR_M1008_s N_VPWR_M1006_s
+ N_VPWR_M1013_d N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_341_n VPWR N_VPWR_c_342_n N_VPWR_c_343_n
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_335_n
+ PM_SKY130_FD_SC_HS__NAND2B_4%VPWR
x_PM_SKY130_FD_SC_HS__NAND2B_4%Y N_Y_M1000_d N_Y_M1010_d N_Y_M1003_d N_Y_M1002_s
+ N_Y_c_400_n N_Y_c_401_n N_Y_c_406_n N_Y_c_412_n N_Y_c_397_n N_Y_c_471_p
+ N_Y_c_416_n N_Y_c_395_n N_Y_c_396_n N_Y_c_433_n N_Y_c_437_n N_Y_c_399_n
+ N_Y_c_424_n Y Y N_Y_c_441_n Y N_Y_c_443_n PM_SKY130_FD_SC_HS__NAND2B_4%Y
x_PM_SKY130_FD_SC_HS__NAND2B_4%VGND N_VGND_M1012_d N_VGND_M1001_s N_VGND_M1009_s
+ N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n VGND
+ N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n
+ N_VGND_c_485_n N_VGND_c_486_n PM_SKY130_FD_SC_HS__NAND2B_4%VGND
x_PM_SKY130_FD_SC_HS__NAND2B_4%A_243_74# N_A_243_74#_M1000_s N_A_243_74#_M1007_s
+ N_A_243_74#_M1014_s N_A_243_74#_M1004_d N_A_243_74#_M1011_d
+ N_A_243_74#_c_545_n N_A_243_74#_c_546_n N_A_243_74#_c_547_n
+ N_A_243_74#_c_560_n N_A_243_74#_c_548_n N_A_243_74#_c_567_n
+ N_A_243_74#_c_575_n N_A_243_74#_c_569_n N_A_243_74#_c_549_n
+ N_A_243_74#_c_550_n N_A_243_74#_c_551_n N_A_243_74#_c_552_n
+ N_A_243_74#_c_553_n PM_SKY130_FD_SC_HS__NAND2B_4%A_243_74#
cc_1 VNB N_A_N_M1012_g 0.0336637f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_2 VNB N_A_N_c_86_n 0.014611f $X=-0.19 $Y=-0.245 $X2=1.53 $Y2=1.65
cc_3 VNB N_A_N_c_87_n 0.030747f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.512
cc_4 VNB N_A_N_c_88_n 0.0181524f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.532
cc_5 VNB N_A_N_c_89_n 0.0379072f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.512
cc_6 VNB N_A_N_c_90_n 0.0146212f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.465
cc_7 VNB N_A_31_74#_c_138_n 0.0163718f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=2.26
cc_8 VNB N_A_31_74#_c_139_n 0.0135187f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.765
cc_9 VNB N_A_31_74#_c_140_n 0.00859217f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.26
cc_10 VNB N_A_31_74#_c_141_n 0.0137758f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.26
cc_11 VNB N_A_31_74#_c_142_n 0.014738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_31_74#_c_143_n 0.0147701f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_13 VNB N_A_31_74#_c_144_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_31_74#_c_145_n 0.0181961f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.54
cc_15 VNB N_A_31_74#_c_146_n 0.00862043f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_16 VNB N_A_31_74#_c_147_n 0.00750487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_31_74#_c_148_n 0.00706303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_31_74#_c_149_n 8.53246e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_31_74#_c_150_n 0.0827825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_M1001_g 0.0199761f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_21 VNB N_B_c_256_n 0.0263567f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.765
cc_22 VNB N_B_c_257_n 0.0139238f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=2.26
cc_23 VNB N_B_M1004_g 0.0212517f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.65
cc_24 VNB N_B_M1009_g 0.0267716f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.512
cc_25 VNB N_B_M1011_g 0.0356645f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.512
cc_26 VNB B 0.0160381f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_27 VNB N_B_c_262_n 0.130318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_263_n 0.00122182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_335_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_395_n 0.00458756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_396_n 0.00491883f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_32 VNB N_VGND_c_476_n 0.0108651f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.26
cc_33 VNB N_VGND_c_477_n 0.00536643f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_34 VNB N_VGND_c_478_n 0.0161561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_479_n 0.0124478f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.465
cc_36 VNB N_VGND_c_480_n 0.0180274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_481_n 0.0626005f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.54
cc_38 VNB N_VGND_c_482_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_483_n 0.326567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_484_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_485_n 0.00612757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_486_n 0.0127911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_243_74#_c_545_n 0.003759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_243_74#_c_546_n 0.00230691f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.512
cc_45 VNB N_A_243_74#_c_547_n 0.00404005f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.465
cc_46 VNB N_A_243_74#_c_548_n 0.00522428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_243_74#_c_549_n 0.00223498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_243_74#_c_550_n 0.0145845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_243_74#_c_551_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_243_74#_c_552_n 0.00203753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_243_74#_c_553_n 0.00230008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_A_N_c_91_n 0.0175905f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.765
cc_53 VPB N_A_N_c_86_n 0.014907f $X=-0.19 $Y=1.66 $X2=1.53 $Y2=1.65
cc_54 VPB N_A_N_c_93_n 0.016184f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.765
cc_55 VPB N_A_N_c_87_n 0.0173099f $X=-0.19 $Y=1.66 $X2=1.08 $Y2=1.512
cc_56 VPB N_A_N_c_88_n 0.00462798f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.532
cc_57 VPB N_A_N_c_89_n 0.0189391f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.512
cc_58 VPB N_A_N_c_90_n 0.0249809f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.465
cc_59 VPB N_A_31_74#_c_151_n 0.019739f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_60 VPB N_A_31_74#_c_152_n 0.0197822f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.465
cc_61 VPB N_A_31_74#_c_153_n 0.00394633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_31_74#_c_148_n 0.00496929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_31_74#_c_155_n 0.00190852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_31_74#_c_150_n 0.0343627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_B_c_264_n 0.0182112f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_66 VPB N_B_c_265_n 0.0181238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB B 0.0129818f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.54
cc_68 VPB N_B_c_262_n 0.0146139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_B_c_263_n 0.00793085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_336_n 0.0757795f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_71 VPB N_VPWR_c_337_n 0.0170951f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.512
cc_72 VPB N_VPWR_c_338_n 0.0127608f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.512
cc_73 VPB N_VPWR_c_339_n 0.0498794f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_74 VPB N_VPWR_c_340_n 0.0208961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_341_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.54
cc_76 VPB N_VPWR_c_342_n 0.0159859f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.54
cc_77 VPB N_VPWR_c_343_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_344_n 0.0119958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_345_n 0.0251007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_346_n 0.0498477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_335_n 0.0858294f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_Y_c_397_n 0.00587584f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.465
cc_83 VPB N_Y_c_396_n 0.00909692f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.54
cc_84 VPB N_Y_c_399_n 0.00290132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 N_A_N_c_86_n N_A_31_74#_c_140_n 0.0115625f $X=1.53 $Y=1.65 $X2=0 $Y2=0
cc_86 N_A_N_c_88_n N_A_31_74#_c_140_n 0.0019215f $X=1.17 $Y=1.532 $X2=0 $Y2=0
cc_87 N_A_N_c_93_n N_A_31_74#_c_151_n 0.0134593f $X=1.62 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_N_M1012_g N_A_31_74#_c_144_n 0.00159319f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A_N_M1012_g N_A_31_74#_c_145_n 0.0146791f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A_N_c_86_n N_A_31_74#_c_145_n 6.14897e-19 $X=1.53 $Y=1.65 $X2=0 $Y2=0
cc_91 N_A_N_c_87_n N_A_31_74#_c_145_n 0.0184042f $X=1.08 $Y=1.512 $X2=0 $Y2=0
cc_92 N_A_N_c_89_n N_A_31_74#_c_145_n 0.00129703f $X=0.59 $Y=1.512 $X2=0 $Y2=0
cc_93 N_A_N_c_90_n N_A_31_74#_c_145_n 0.0558012f $X=0.95 $Y=1.465 $X2=0 $Y2=0
cc_94 N_A_N_c_89_n N_A_31_74#_c_146_n 0.00612466f $X=0.59 $Y=1.512 $X2=0 $Y2=0
cc_95 N_A_N_c_90_n N_A_31_74#_c_146_n 0.0216392f $X=0.95 $Y=1.465 $X2=0 $Y2=0
cc_96 N_A_N_c_91_n N_A_31_74#_c_153_n 0.00896608f $X=1.17 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A_N_c_86_n N_A_31_74#_c_153_n 0.00131774f $X=1.53 $Y=1.65 $X2=0 $Y2=0
cc_98 N_A_N_c_93_n N_A_31_74#_c_153_n 0.00885631f $X=1.62 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_N_M1012_g N_A_31_74#_c_147_n 0.00337332f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_N_c_88_n N_A_31_74#_c_147_n 0.00328335f $X=1.17 $Y=1.532 $X2=0 $Y2=0
cc_101 N_A_N_c_90_n N_A_31_74#_c_147_n 0.0102699f $X=0.95 $Y=1.465 $X2=0 $Y2=0
cc_102 N_A_N_c_86_n N_A_31_74#_c_148_n 0.0139508f $X=1.53 $Y=1.65 $X2=0 $Y2=0
cc_103 N_A_N_c_91_n N_A_31_74#_c_155_n 0.00194928f $X=1.17 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_N_c_86_n N_A_31_74#_c_155_n 0.0070871f $X=1.53 $Y=1.65 $X2=0 $Y2=0
cc_105 N_A_N_c_93_n N_A_31_74#_c_155_n 0.00268655f $X=1.62 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A_N_c_88_n N_A_31_74#_c_155_n 2.98825e-19 $X=1.17 $Y=1.532 $X2=0 $Y2=0
cc_107 N_A_N_c_90_n N_A_31_74#_c_155_n 0.00766656f $X=0.95 $Y=1.465 $X2=0 $Y2=0
cc_108 N_A_N_c_86_n N_A_31_74#_c_149_n 0.00716973f $X=1.53 $Y=1.65 $X2=0 $Y2=0
cc_109 N_A_N_c_88_n N_A_31_74#_c_149_n 0.00470418f $X=1.17 $Y=1.532 $X2=0 $Y2=0
cc_110 N_A_N_c_90_n N_A_31_74#_c_149_n 0.0218137f $X=0.95 $Y=1.465 $X2=0 $Y2=0
cc_111 N_A_N_c_86_n N_A_31_74#_c_150_n 0.00696242f $X=1.53 $Y=1.65 $X2=0 $Y2=0
cc_112 N_A_N_c_91_n N_VPWR_c_336_n 0.0061881f $X=1.17 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_N_c_89_n N_VPWR_c_336_n 0.00418355f $X=0.59 $Y=1.512 $X2=0 $Y2=0
cc_114 N_A_N_c_90_n N_VPWR_c_336_n 0.054616f $X=0.95 $Y=1.465 $X2=0 $Y2=0
cc_115 N_A_N_c_93_n N_VPWR_c_337_n 0.0109593f $X=1.62 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_N_c_91_n N_VPWR_c_340_n 0.00393873f $X=1.17 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_N_c_93_n N_VPWR_c_340_n 0.00393873f $X=1.62 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A_N_c_91_n N_VPWR_c_335_n 0.00462577f $X=1.17 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_N_c_93_n N_VPWR_c_335_n 0.00462577f $X=1.62 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_N_M1012_g N_VGND_c_476_n 0.013544f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_N_M1012_g N_VGND_c_480_n 0.00383152f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A_N_M1012_g N_VGND_c_483_n 0.00761264f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_N_M1012_g N_A_243_74#_c_545_n 7.29222e-19 $X=0.515 $Y=0.74 $X2=0
+ $Y2=0
cc_124 N_A_N_M1012_g N_A_243_74#_c_547_n 6.35506e-19 $X=0.515 $Y=0.74 $X2=0
+ $Y2=0
cc_125 N_A_31_74#_c_143_n N_B_M1001_g 0.0166524f $X=3 $Y=1.185 $X2=0 $Y2=0
cc_126 N_A_31_74#_c_148_n N_B_c_257_n 2.22559e-19 $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A_31_74#_c_150_n N_B_c_257_n 0.0166524f $X=2.985 $Y=1.475 $X2=0 $Y2=0
cc_128 N_A_31_74#_c_153_n N_VPWR_c_336_n 0.0289748f $X=1.395 $Y=2.115 $X2=0
+ $Y2=0
cc_129 N_A_31_74#_c_151_n N_VPWR_c_337_n 0.01919f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_31_74#_c_153_n N_VPWR_c_337_n 0.0504069f $X=1.395 $Y=2.115 $X2=0
+ $Y2=0
cc_131 N_A_31_74#_c_148_n N_VPWR_c_337_n 0.0251163f $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A_31_74#_c_155_n N_VPWR_c_337_n 0.00488691f $X=1.395 $Y=1.95 $X2=0
+ $Y2=0
cc_133 N_A_31_74#_c_153_n N_VPWR_c_340_n 0.00664674f $X=1.395 $Y=2.115 $X2=0
+ $Y2=0
cc_134 N_A_31_74#_c_151_n N_VPWR_c_345_n 0.00413917f $X=2.155 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_31_74#_c_152_n N_VPWR_c_345_n 0.00413917f $X=2.985 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_31_74#_c_152_n N_VPWR_c_346_n 0.0156712f $X=2.985 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_31_74#_c_151_n N_VPWR_c_335_n 0.00820334f $X=2.155 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_31_74#_c_152_n N_VPWR_c_335_n 0.00815719f $X=2.985 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_31_74#_c_153_n N_VPWR_c_335_n 0.00995652f $X=1.395 $Y=2.115 $X2=0
+ $Y2=0
cc_140 N_A_31_74#_c_138_n N_Y_c_400_n 0.011255f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A_31_74#_c_139_n N_Y_c_401_n 6.06204e-19 $X=1.93 $Y=1.26 $X2=0 $Y2=0
cc_142 N_A_31_74#_c_141_n N_Y_c_401_n 0.00745896f $X=2.005 $Y=1.185 $X2=0 $Y2=0
cc_143 N_A_31_74#_c_142_n N_Y_c_401_n 0.00784525f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_144 N_A_31_74#_c_148_n N_Y_c_401_n 0.0474062f $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A_31_74#_c_150_n N_Y_c_401_n 0.0136143f $X=2.985 $Y=1.475 $X2=0 $Y2=0
cc_146 N_A_31_74#_c_138_n N_Y_c_406_n 0.00213594f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_147 N_A_31_74#_c_139_n N_Y_c_406_n 0.00555852f $X=1.93 $Y=1.26 $X2=0 $Y2=0
cc_148 N_A_31_74#_c_140_n N_Y_c_406_n 9.64687e-19 $X=1.65 $Y=1.26 $X2=0 $Y2=0
cc_149 N_A_31_74#_c_145_n N_Y_c_406_n 0.00258252f $X=1.285 $Y=1.045 $X2=0 $Y2=0
cc_150 N_A_31_74#_c_147_n N_Y_c_406_n 0.0103078f $X=1.37 $Y=1.43 $X2=0 $Y2=0
cc_151 N_A_31_74#_c_148_n N_Y_c_406_n 0.0211885f $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A_31_74#_c_148_n N_Y_c_412_n 0.0474415f $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A_31_74#_c_150_n N_Y_c_412_n 0.0160066f $X=2.985 $Y=1.475 $X2=0 $Y2=0
cc_154 N_A_31_74#_c_151_n N_Y_c_397_n 4.34144e-19 $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_31_74#_c_152_n N_Y_c_397_n 4.33747e-19 $X=2.985 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A_31_74#_c_152_n N_Y_c_416_n 0.0199901f $X=2.985 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_31_74#_c_148_n N_Y_c_416_n 0.0127017f $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A_31_74#_c_143_n N_Y_c_395_n 0.00783312f $X=3 $Y=1.185 $X2=0 $Y2=0
cc_159 N_A_31_74#_c_148_n N_Y_c_395_n 0.0135868f $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A_31_74#_c_150_n N_Y_c_395_n 0.00489222f $X=2.985 $Y=1.475 $X2=0 $Y2=0
cc_161 N_A_31_74#_c_152_n N_Y_c_396_n 0.0029796f $X=2.985 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_31_74#_c_148_n N_Y_c_396_n 0.0178989f $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A_31_74#_c_150_n N_Y_c_396_n 0.00839068f $X=2.985 $Y=1.475 $X2=0 $Y2=0
cc_164 N_A_31_74#_c_148_n N_Y_c_424_n 0.0252592f $X=2.91 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A_31_74#_c_150_n N_Y_c_424_n 0.0122905f $X=2.985 $Y=1.475 $X2=0 $Y2=0
cc_166 N_A_31_74#_c_145_n N_VGND_M1012_d 0.00328964f $X=1.285 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_167 N_A_31_74#_c_138_n N_VGND_c_476_n 8.77482e-19 $X=1.575 $Y=1.185 $X2=0
+ $Y2=0
cc_168 N_A_31_74#_c_144_n N_VGND_c_476_n 0.0164982f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_169 N_A_31_74#_c_145_n N_VGND_c_476_n 0.0219827f $X=1.285 $Y=1.045 $X2=0
+ $Y2=0
cc_170 N_A_31_74#_c_144_n N_VGND_c_480_n 0.011066f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_171 N_A_31_74#_c_138_n N_VGND_c_481_n 0.00278271f $X=1.575 $Y=1.185 $X2=0
+ $Y2=0
cc_172 N_A_31_74#_c_141_n N_VGND_c_481_n 0.00278247f $X=2.005 $Y=1.185 $X2=0
+ $Y2=0
cc_173 N_A_31_74#_c_142_n N_VGND_c_481_n 0.00278247f $X=2.435 $Y=1.185 $X2=0
+ $Y2=0
cc_174 N_A_31_74#_c_143_n N_VGND_c_481_n 0.00278247f $X=3 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A_31_74#_c_138_n N_VGND_c_483_n 0.00358427f $X=1.575 $Y=1.185 $X2=0
+ $Y2=0
cc_176 N_A_31_74#_c_141_n N_VGND_c_483_n 0.00353427f $X=2.005 $Y=1.185 $X2=0
+ $Y2=0
cc_177 N_A_31_74#_c_142_n N_VGND_c_483_n 0.00354622f $X=2.435 $Y=1.185 $X2=0
+ $Y2=0
cc_178 N_A_31_74#_c_143_n N_VGND_c_483_n 0.00354719f $X=3 $Y=1.185 $X2=0 $Y2=0
cc_179 N_A_31_74#_c_144_n N_VGND_c_483_n 0.00915947f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_180 N_A_31_74#_c_145_n N_A_243_74#_M1000_s 0.00436281f $X=1.285 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_181 N_A_31_74#_c_145_n N_A_243_74#_c_545_n 0.0211188f $X=1.285 $Y=1.045 $X2=0
+ $Y2=0
cc_182 N_A_31_74#_c_138_n N_A_243_74#_c_546_n 0.013422f $X=1.575 $Y=1.185 $X2=0
+ $Y2=0
cc_183 N_A_31_74#_c_141_n N_A_243_74#_c_546_n 0.00815411f $X=2.005 $Y=1.185
+ $X2=0 $Y2=0
cc_184 N_A_31_74#_c_138_n N_A_243_74#_c_560_n 6.13499e-19 $X=1.575 $Y=1.185
+ $X2=0 $Y2=0
cc_185 N_A_31_74#_c_141_n N_A_243_74#_c_560_n 0.00708959f $X=2.005 $Y=1.185
+ $X2=0 $Y2=0
cc_186 N_A_31_74#_c_142_n N_A_243_74#_c_560_n 0.00750562f $X=2.435 $Y=1.185
+ $X2=0 $Y2=0
cc_187 N_A_31_74#_c_143_n N_A_243_74#_c_560_n 7.13474e-19 $X=3 $Y=1.185 $X2=0
+ $Y2=0
cc_188 N_A_31_74#_c_150_n N_A_243_74#_c_560_n 6.12873e-19 $X=2.985 $Y=1.475
+ $X2=0 $Y2=0
cc_189 N_A_31_74#_c_142_n N_A_243_74#_c_548_n 0.00885191f $X=2.435 $Y=1.185
+ $X2=0 $Y2=0
cc_190 N_A_31_74#_c_143_n N_A_243_74#_c_548_n 0.0107003f $X=3 $Y=1.185 $X2=0
+ $Y2=0
cc_191 N_A_31_74#_c_142_n N_A_243_74#_c_567_n 6.79059e-19 $X=2.435 $Y=1.185
+ $X2=0 $Y2=0
cc_192 N_A_31_74#_c_143_n N_A_243_74#_c_567_n 0.00540996f $X=3 $Y=1.185 $X2=0
+ $Y2=0
cc_193 N_A_31_74#_c_143_n N_A_243_74#_c_569_n 0.00210741f $X=3 $Y=1.185 $X2=0
+ $Y2=0
cc_194 N_A_31_74#_c_141_n N_A_243_74#_c_552_n 0.00187501f $X=2.005 $Y=1.185
+ $X2=0 $Y2=0
cc_195 N_A_31_74#_c_142_n N_A_243_74#_c_552_n 0.00187501f $X=2.435 $Y=1.185
+ $X2=0 $Y2=0
cc_196 N_B_c_265_n N_VPWR_c_339_n 0.00371973f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_197 B N_VPWR_c_339_n 0.0243138f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_198 N_B_c_262_n N_VPWR_c_339_n 0.00116212f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_199 N_B_c_264_n N_VPWR_c_343_n 0.00461464f $X=4.735 $Y=1.765 $X2=0 $Y2=0
cc_200 N_B_c_265_n N_VPWR_c_343_n 0.00445602f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_201 N_B_c_256_n N_VPWR_c_346_n 9.72602e-19 $X=3.855 $Y=1.465 $X2=0 $Y2=0
cc_202 N_B_c_257_n N_VPWR_c_346_n 8.52878e-19 $X=3.505 $Y=1.465 $X2=0 $Y2=0
cc_203 N_B_c_264_n N_VPWR_c_346_n 0.0045193f $X=4.735 $Y=1.765 $X2=0 $Y2=0
cc_204 N_B_c_264_n N_VPWR_c_335_n 0.009128f $X=4.735 $Y=1.765 $X2=0 $Y2=0
cc_205 N_B_c_265_n N_VPWR_c_335_n 0.00860756f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_206 N_B_M1001_g N_Y_c_395_n 0.00807839f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B_M1004_g N_Y_c_395_n 0.00390557f $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B_M1001_g N_Y_c_396_n 0.00107252f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B_c_256_n N_Y_c_396_n 0.0139602f $X=3.855 $Y=1.465 $X2=0 $Y2=0
cc_210 N_B_c_257_n N_Y_c_396_n 0.00977419f $X=3.505 $Y=1.465 $X2=0 $Y2=0
cc_211 N_B_M1004_g N_Y_c_396_n 9.32683e-19 $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B_c_288_p N_Y_c_396_n 0.0241378f $X=4.445 $Y=1.54 $X2=0 $Y2=0
cc_213 N_B_c_264_n N_Y_c_433_n 0.0163174f $X=4.735 $Y=1.765 $X2=0 $Y2=0
cc_214 N_B_c_262_n N_Y_c_433_n 0.00681852f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_215 N_B_c_263_n N_Y_c_433_n 0.0267106f $X=4.925 $Y=1.54 $X2=0 $Y2=0
cc_216 N_B_c_288_p N_Y_c_433_n 0.0114511f $X=4.445 $Y=1.54 $X2=0 $Y2=0
cc_217 N_B_c_265_n N_Y_c_437_n 0.00220431f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_218 N_B_c_262_n N_Y_c_437_n 0.00142563f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_219 N_B_c_263_n N_Y_c_437_n 0.024327f $X=4.925 $Y=1.54 $X2=0 $Y2=0
cc_220 N_B_c_265_n N_Y_c_399_n 0.0086185f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_221 N_B_c_256_n N_Y_c_441_n 0.00805051f $X=3.855 $Y=1.465 $X2=0 $Y2=0
cc_222 N_B_c_288_p N_Y_c_441_n 0.0220598f $X=4.445 $Y=1.54 $X2=0 $Y2=0
cc_223 N_B_c_264_n N_Y_c_443_n 0.0029836f $X=4.735 $Y=1.765 $X2=0 $Y2=0
cc_224 N_B_c_262_n N_Y_c_443_n 0.00805051f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_225 N_B_M1001_g N_VGND_c_477_n 0.00246766f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B_M1004_g N_VGND_c_477_n 0.00655891f $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B_M1009_g N_VGND_c_477_n 3.63592e-19 $X=4.36 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B_M1004_g N_VGND_c_478_n 0.00281948f $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B_M1009_g N_VGND_c_478_n 0.00433834f $X=4.36 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B_M1009_g N_VGND_c_479_n 0.00482335f $X=4.36 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B_M1011_g N_VGND_c_479_n 0.00669543f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B_M1001_g N_VGND_c_481_n 0.00328073f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_233 N_B_M1011_g N_VGND_c_482_n 0.00434272f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B_M1001_g N_VGND_c_483_n 0.00426855f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B_M1004_g N_VGND_c_483_n 0.00363526f $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B_M1009_g N_VGND_c_483_n 0.00824753f $X=4.36 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B_M1011_g N_VGND_c_483_n 0.00828717f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B_M1001_g N_A_243_74#_c_548_n 0.00320891f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B_M1001_g N_A_243_74#_c_567_n 0.00494934f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B_M1004_g N_A_243_74#_c_567_n 2.75259e-19 $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B_M1001_g N_A_243_74#_c_575_n 0.00915554f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_242 N_B_c_256_n N_A_243_74#_c_575_n 0.00357964f $X=3.855 $Y=1.465 $X2=0 $Y2=0
cc_243 N_B_M1004_g N_A_243_74#_c_575_n 0.0108383f $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_244 N_B_c_288_p N_A_243_74#_c_575_n 0.00485175f $X=4.445 $Y=1.54 $X2=0 $Y2=0
cc_245 N_B_M1001_g N_A_243_74#_c_569_n 7.30706e-19 $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_246 N_B_M1004_g N_A_243_74#_c_549_n 5.30282e-19 $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_247 N_B_M1009_g N_A_243_74#_c_549_n 0.00555458f $X=4.36 $Y=0.74 $X2=0 $Y2=0
cc_248 N_B_M1009_g N_A_243_74#_c_550_n 0.0142398f $X=4.36 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B_M1011_g N_A_243_74#_c_550_n 0.0143229f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_250 B N_A_243_74#_c_550_n 0.0289285f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B_c_262_n N_A_243_74#_c_550_n 0.0180748f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_252 N_B_c_288_p N_A_243_74#_c_550_n 0.0764136f $X=4.445 $Y=1.54 $X2=0 $Y2=0
cc_253 N_B_M1011_g N_A_243_74#_c_551_n 0.0138506f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_254 N_B_M1001_g N_A_243_74#_c_553_n 9.2198e-19 $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B_M1004_g N_A_243_74#_c_553_n 0.00584308f $X=3.93 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B_M1009_g N_A_243_74#_c_553_n 0.00930967f $X=4.36 $Y=0.74 $X2=0 $Y2=0
cc_257 N_B_c_262_n N_A_243_74#_c_553_n 0.00232957f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_258 N_B_c_288_p N_A_243_74#_c_553_n 0.0271869f $X=4.445 $Y=1.54 $X2=0 $Y2=0
cc_259 N_VPWR_c_337_n N_Y_c_397_n 0.0320109f $X=1.93 $Y=2.015 $X2=0 $Y2=0
cc_260 N_VPWR_c_345_n N_Y_c_397_n 0.0271295f $X=3.045 $Y=2.867 $X2=0 $Y2=0
cc_261 N_VPWR_c_346_n N_Y_c_397_n 0.0286308f $X=4.645 $Y=2.867 $X2=0 $Y2=0
cc_262 N_VPWR_c_335_n N_Y_c_397_n 0.0224555f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_263 N_VPWR_M1006_s N_Y_c_416_n 0.00562147f $X=3.06 $Y=1.84 $X2=0 $Y2=0
cc_264 N_VPWR_c_346_n N_Y_c_416_n 0.0152517f $X=4.645 $Y=2.867 $X2=0 $Y2=0
cc_265 N_VPWR_M1006_s N_Y_c_396_n 6.79886e-19 $X=3.06 $Y=1.84 $X2=0 $Y2=0
cc_266 N_VPWR_M1006_s N_Y_c_433_n 0.011768f $X=3.06 $Y=1.84 $X2=0 $Y2=0
cc_267 N_VPWR_c_339_n N_Y_c_399_n 0.0318792f $X=5.435 $Y=2.115 $X2=0 $Y2=0
cc_268 N_VPWR_c_343_n N_Y_c_399_n 0.0145938f $X=5.315 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_c_346_n N_Y_c_399_n 0.00167954f $X=4.645 $Y=2.867 $X2=0 $Y2=0
cc_270 N_VPWR_c_335_n N_Y_c_399_n 0.0120466f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_271 N_VPWR_M1006_s Y 0.0102263f $X=3.06 $Y=1.84 $X2=0 $Y2=0
cc_272 N_VPWR_c_346_n Y 0.0331229f $X=4.645 $Y=2.867 $X2=0 $Y2=0
cc_273 N_VPWR_M1006_s N_Y_c_441_n 0.0149516f $X=3.06 $Y=1.84 $X2=0 $Y2=0
cc_274 N_VPWR_c_346_n N_Y_c_441_n 0.0787788f $X=4.645 $Y=2.867 $X2=0 $Y2=0
cc_275 N_VPWR_M1006_s N_Y_c_443_n 0.00728674f $X=3.06 $Y=1.84 $X2=0 $Y2=0
cc_276 N_Y_c_395_n N_VGND_M1001_s 0.00126218f $X=3.285 $Y=1.175 $X2=0 $Y2=0
cc_277 N_Y_c_401_n N_A_243_74#_M1007_s 0.00176461f $X=2.555 $Y=1.175 $X2=0 $Y2=0
cc_278 N_Y_c_395_n N_A_243_74#_M1014_s 0.00175965f $X=3.285 $Y=1.175 $X2=0 $Y2=0
cc_279 N_Y_M1000_d N_A_243_74#_c_546_n 0.00193374f $X=1.65 $Y=0.37 $X2=0 $Y2=0
cc_280 N_Y_c_400_n N_A_243_74#_c_546_n 0.0118362f $X=1.79 $Y=0.82 $X2=0 $Y2=0
cc_281 N_Y_c_401_n N_A_243_74#_c_546_n 0.00270072f $X=2.555 $Y=1.175 $X2=0 $Y2=0
cc_282 N_Y_c_401_n N_A_243_74#_c_560_n 0.0170464f $X=2.555 $Y=1.175 $X2=0 $Y2=0
cc_283 N_Y_M1010_d N_A_243_74#_c_548_n 0.00367075f $X=2.51 $Y=0.37 $X2=0 $Y2=0
cc_284 N_Y_c_401_n N_A_243_74#_c_548_n 0.00270072f $X=2.555 $Y=1.175 $X2=0 $Y2=0
cc_285 N_Y_c_471_p N_A_243_74#_c_548_n 0.0189799f $X=2.725 $Y=0.82 $X2=0 $Y2=0
cc_286 N_Y_c_395_n N_A_243_74#_c_548_n 0.00270072f $X=3.285 $Y=1.175 $X2=0 $Y2=0
cc_287 N_Y_c_395_n N_A_243_74#_c_575_n 0.0170542f $X=3.285 $Y=1.175 $X2=0 $Y2=0
cc_288 N_Y_c_395_n N_A_243_74#_c_569_n 0.0174882f $X=3.285 $Y=1.175 $X2=0 $Y2=0
cc_289 N_Y_c_395_n N_A_243_74#_c_553_n 0.00204498f $X=3.285 $Y=1.175 $X2=0 $Y2=0
cc_290 N_VGND_c_476_n N_A_243_74#_c_545_n 0.020109f $X=0.73 $Y=0.57 $X2=0 $Y2=0
cc_291 N_VGND_c_481_n N_A_243_74#_c_546_n 0.0377951f $X=3.55 $Y=0 $X2=0 $Y2=0
cc_292 N_VGND_c_483_n N_A_243_74#_c_546_n 0.0212998f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_293 N_VGND_c_476_n N_A_243_74#_c_547_n 0.0101239f $X=0.73 $Y=0.57 $X2=0 $Y2=0
cc_294 N_VGND_c_481_n N_A_243_74#_c_547_n 0.0183077f $X=3.55 $Y=0 $X2=0 $Y2=0
cc_295 N_VGND_c_483_n N_A_243_74#_c_547_n 0.0100461f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_296 N_VGND_c_477_n N_A_243_74#_c_548_n 0.011924f $X=3.715 $Y=0.495 $X2=0
+ $Y2=0
cc_297 N_VGND_c_481_n N_A_243_74#_c_548_n 0.0654994f $X=3.55 $Y=0 $X2=0 $Y2=0
cc_298 N_VGND_c_483_n N_A_243_74#_c_548_n 0.0364513f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_299 N_VGND_M1001_s N_A_243_74#_c_575_n 0.00611887f $X=3.505 $Y=0.37 $X2=0
+ $Y2=0
cc_300 N_VGND_c_477_n N_A_243_74#_c_575_n 0.0203034f $X=3.715 $Y=0.495 $X2=0
+ $Y2=0
cc_301 N_VGND_c_478_n N_A_243_74#_c_575_n 0.00125985f $X=4.48 $Y=0 $X2=0 $Y2=0
cc_302 N_VGND_c_481_n N_A_243_74#_c_575_n 0.00189877f $X=3.55 $Y=0 $X2=0 $Y2=0
cc_303 N_VGND_c_483_n N_A_243_74#_c_575_n 0.00719631f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_477_n N_A_243_74#_c_549_n 0.0109457f $X=3.715 $Y=0.495 $X2=0
+ $Y2=0
cc_305 N_VGND_c_478_n N_A_243_74#_c_549_n 0.0124403f $X=4.48 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_479_n N_A_243_74#_c_549_n 0.0184625f $X=5.05 $Y=0.625 $X2=0
+ $Y2=0
cc_307 N_VGND_c_483_n N_A_243_74#_c_549_n 0.00952716f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_308 N_VGND_M1009_s N_A_243_74#_c_550_n 0.0100716f $X=4.435 $Y=0.37 $X2=0
+ $Y2=0
cc_309 N_VGND_c_479_n N_A_243_74#_c_550_n 0.0521508f $X=5.05 $Y=0.625 $X2=0
+ $Y2=0
cc_310 N_VGND_c_479_n N_A_243_74#_c_551_n 0.0173886f $X=5.05 $Y=0.625 $X2=0
+ $Y2=0
cc_311 N_VGND_c_482_n N_A_243_74#_c_551_n 0.0145639f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_483_n N_A_243_74#_c_551_n 0.0119984f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_c_481_n N_A_243_74#_c_552_n 0.0234416f $X=3.55 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_483_n N_A_243_74#_c_552_n 0.0125934f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_478_n N_A_243_74#_c_553_n 6.44141e-19 $X=4.48 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_c_483_n N_A_243_74#_c_553_n 0.00173608f $X=5.52 $Y=0 $X2=0 $Y2=0
