* File: sky130_fd_sc_hs__a311oi_1.spice
* Created: Thu Aug 27 20:28:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a311oi_1.pex.spice"
.subckt sky130_fd_sc_hs__a311oi_1  VNB VPB A3 A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1004 A_159_74# N_A3_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75002.2
+ A=0.111 P=1.78 MULT=1
MM1002 A_231_74# N_A2_M1002_g A_159_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.0777 PD=1.13 PS=0.95 NRD=22.692 NRS=8.1 M=1 R=4.93333 SA=75000.6
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1006_d N_A1_M1006_g A_231_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.1443 PD=1.13 PS=1.13 NRD=3.24 NRS=22.692 M=1 R=4.93333 SA=75001.1
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_B1_M1009_g N_Y_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=3.24 NRS=14.592 M=1 R=4.93333
+ SA=75001.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75002.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_156_368#_M1000_d N_A3_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_156_368#_M1000_d VPB PSHORT L=0.15 W=1.12
+ AD=0.2688 AS=0.168 PD=1.6 PS=1.42 NRD=17.5724 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1007 N_A_156_368#_M1007_d N_A1_M1007_g N_VPWR_M1001_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2688 PD=1.42 PS=1.6 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75001.3 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1008 A_462_368# N_B1_M1008_g N_A_156_368#_M1007_d VPB PSHORT L=0.15 W=1.12
+ AD=0.1848 AS=0.168 PD=1.45 PS=1.42 NRD=19.3454 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1005_d N_C1_M1005_g A_462_368# VPB PSHORT L=0.15 W=1.12 AD=0.308
+ AS=0.1848 PD=2.79 PS=1.45 NRD=1.7533 NRS=19.3454 M=1 R=7.46667 SA=75002.2
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__a311oi_1.pxi.spice"
*
.ends
*
*
