* File: sky130_fd_sc_hs__bufbuf_8.pex.spice
* Created: Tue Sep  1 19:57:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__BUFBUF_8%A 3 5 7 8 12
c34 5 0 1.95957e-19 $X=0.505 $Y=1.765
c35 3 0 8.22433e-20 $X=0.495 $Y=0.835
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.515 $X2=0.405 $Y2=1.515
r37 8 12 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.405 $Y2=1.565
r38 5 11 52.4131 $w=2.96e-07 $l=2.93684e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.41 $Y2=1.515
r39 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
r40 1 11 38.5718 $w=2.96e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.41 $Y2=1.515
r41 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__BUFBUF_8%A_27_112# 1 2 7 9 12 16 18 20 22 24 25 26
+ 27
r71 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.465 $X2=0.975 $Y2=1.465
r72 26 32 9.02499 $w=2.87e-07 $l=2.13014e-07 $layer=LI1_cond $X=0.835 $Y=1.63
+ $X2=0.945 $Y2=1.465
r73 26 27 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.835 $Y=1.63
+ $X2=0.835 $Y2=1.95
r74 24 32 15.7282 $w=2.87e-07 $l=4.5722e-07 $layer=LI1_cond $X=0.75 $Y=1.095
+ $X2=0.945 $Y2=1.465
r75 24 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.75 $Y=1.095
+ $X2=0.445 $Y2=1.095
r76 23 29 3.51781 $w=2.5e-07 $l=1.33e-07 $layer=LI1_cond $X=0.38 $Y=2.075
+ $X2=0.247 $Y2=2.075
r77 22 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.75 $Y=2.075
+ $X2=0.835 $Y2=1.95
r78 22 23 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=2.075
+ $X2=0.38 $Y2=2.075
r79 18 29 3.30621 $w=2.65e-07 $l=1.25e-07 $layer=LI1_cond $X=0.247 $Y=2.2
+ $X2=0.247 $Y2=2.075
r80 18 20 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=0.247 $Y=2.2
+ $X2=0.247 $Y2=2.535
r81 14 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r82 14 16 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.835
r83 10 33 38.5916 $w=2.93e-07 $l=2.07123e-07 $layer=POLY_cond $X=1.075 $Y=1.3
+ $X2=0.98 $Y2=1.465
r84 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.075 $Y=1.3
+ $X2=1.075 $Y2=0.74
r85 7 33 60.7998 $w=2.93e-07 $l=3.24037e-07 $layer=POLY_cond $X=1.03 $Y=1.765
+ $X2=0.98 $Y2=1.465
r86 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.03 $Y=1.765
+ $X2=1.03 $Y2=2.4
r87 2 29 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.06
r88 2 20 600 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.535
r89 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__BUFBUF_8%A_221_368# 1 2 7 9 12 14 16 19 23 25 27 30
+ 34 37 45 49 50 51 52 53 61
c99 51 0 8.22433e-20 $X=1.302 $Y=1.13
c100 49 0 1.95957e-19 $X=1.255 $Y=1.985
c101 23 0 2.25722e-20 $X=2.925 $Y=0.74
r102 61 62 1.82116 $w=3.97e-07 $l=1.5e-08 $layer=POLY_cond $X=2.925 $Y=1.532
+ $X2=2.94 $Y2=1.532
r103 60 61 52.2066 $w=3.97e-07 $l=4.3e-07 $layer=POLY_cond $X=2.495 $Y=1.532
+ $X2=2.925 $Y2=1.532
r104 59 60 0.607053 $w=3.97e-07 $l=5e-09 $layer=POLY_cond $X=2.49 $Y=1.532
+ $X2=2.495 $Y2=1.532
r105 56 57 3.03526 $w=3.97e-07 $l=2.5e-08 $layer=POLY_cond $X=2.04 $Y=1.532
+ $X2=2.065 $Y2=1.532
r106 53 56 12.4421 $w=3.97e-07 $l=1.1887e-07 $layer=POLY_cond $X=1.95 $Y=1.465
+ $X2=2.04 $Y2=1.532
r107 49 50 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=1.985
+ $X2=1.285 $Y2=1.82
r108 46 59 14.5693 $w=3.97e-07 $l=1.2e-07 $layer=POLY_cond $X=2.37 $Y=1.532
+ $X2=2.49 $Y2=1.532
r109 46 57 37.0302 $w=3.97e-07 $l=3.05e-07 $layer=POLY_cond $X=2.37 $Y=1.532
+ $X2=2.065 $Y2=1.532
r110 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.465 $X2=2.37 $Y2=1.465
r111 43 53 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.69 $Y=1.465
+ $X2=1.95 $Y2=1.465
r112 42 45 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.69 $Y=1.465
+ $X2=2.37 $Y2=1.465
r113 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.465 $X2=1.69 $Y2=1.465
r114 40 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=1.465
+ $X2=1.395 $Y2=1.465
r115 40 42 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.48 $Y=1.465
+ $X2=1.69 $Y2=1.465
r116 38 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=1.63
+ $X2=1.395 $Y2=1.465
r117 38 50 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.395 $Y=1.63
+ $X2=1.395 $Y2=1.82
r118 37 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=1.3
+ $X2=1.395 $Y2=1.465
r119 37 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.395 $Y=1.3
+ $X2=1.395 $Y2=1.13
r120 32 51 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=1.302 $Y=0.953
+ $X2=1.302 $Y2=1.13
r121 32 34 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=1.302 $Y=0.953
+ $X2=1.302 $Y2=0.515
r122 28 49 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=1.285 $Y=2.015
+ $X2=1.285 $Y2=1.985
r123 28 30 23.6399 $w=3.88e-07 $l=8e-07 $layer=LI1_cond $X=1.285 $Y=2.015
+ $X2=1.285 $Y2=2.815
r124 25 62 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.94 $Y=1.765
+ $X2=2.94 $Y2=1.532
r125 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.94 $Y=1.765
+ $X2=2.94 $Y2=2.4
r126 21 61 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.925 $Y=1.3
+ $X2=2.925 $Y2=1.532
r127 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.925 $Y=1.3
+ $X2=2.925 $Y2=0.74
r128 17 60 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.495 $Y=1.3
+ $X2=2.495 $Y2=1.532
r129 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.495 $Y=1.3
+ $X2=2.495 $Y2=0.74
r130 14 59 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.49 $Y=1.765
+ $X2=2.49 $Y2=1.532
r131 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.49 $Y=1.765
+ $X2=2.49 $Y2=2.4
r132 10 57 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.065 $Y=1.3
+ $X2=2.065 $Y2=1.532
r133 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.065 $Y=1.3
+ $X2=2.065 $Y2=0.74
r134 7 56 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.04 $Y=1.765
+ $X2=2.04 $Y2=1.532
r135 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.04 $Y=1.765
+ $X2=2.04 $Y2=2.4
r136 2 49 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.84 $X2=1.255 $Y2=1.985
r137 2 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.84 $X2=1.255 $Y2=2.815
r138 1 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.15
+ $Y=0.37 $X2=1.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFBUF_8%A_334_368# 1 2 3 4 15 17 19 22 24 26 29 31
+ 33 36 38 40 43 45 47 50 52 54 55 57 60 64 66 68 69 71 73 75 79 83 86 92 100
+ 102 122
c196 102 0 2.25722e-20 $X=2.71 $Y=0.965
r197 122 123 1.24548 $w=3.87e-07 $l=1e-08 $layer=POLY_cond $X=6.635 $Y=1.532
+ $X2=6.645 $Y2=1.532
r198 121 122 53.5556 $w=3.87e-07 $l=4.3e-07 $layer=POLY_cond $X=6.205 $Y=1.532
+ $X2=6.635 $Y2=1.532
r199 120 121 1.24548 $w=3.87e-07 $l=1e-08 $layer=POLY_cond $X=6.195 $Y=1.532
+ $X2=6.205 $Y2=1.532
r200 117 118 4.98191 $w=3.87e-07 $l=4e-08 $layer=POLY_cond $X=5.705 $Y=1.532
+ $X2=5.745 $Y2=1.532
r201 116 117 51.0646 $w=3.87e-07 $l=4.1e-07 $layer=POLY_cond $X=5.295 $Y=1.532
+ $X2=5.705 $Y2=1.532
r202 115 116 9.96382 $w=3.87e-07 $l=8e-08 $layer=POLY_cond $X=5.215 $Y=1.532
+ $X2=5.295 $Y2=1.532
r203 114 115 46.7054 $w=3.87e-07 $l=3.75e-07 $layer=POLY_cond $X=4.84 $Y=1.532
+ $X2=5.215 $Y2=1.532
r204 113 114 6.85013 $w=3.87e-07 $l=5.5e-08 $layer=POLY_cond $X=4.785 $Y=1.532
+ $X2=4.84 $Y2=1.532
r205 112 113 49.1964 $w=3.87e-07 $l=3.95e-07 $layer=POLY_cond $X=4.39 $Y=1.532
+ $X2=4.785 $Y2=1.532
r206 111 112 4.35917 $w=3.87e-07 $l=3.5e-08 $layer=POLY_cond $X=4.355 $Y=1.532
+ $X2=4.39 $Y2=1.532
r207 110 111 51.6873 $w=3.87e-07 $l=4.15e-07 $layer=POLY_cond $X=3.94 $Y=1.532
+ $X2=4.355 $Y2=1.532
r208 109 110 10.5866 $w=3.87e-07 $l=8.5e-08 $layer=POLY_cond $X=3.855 $Y=1.532
+ $X2=3.94 $Y2=1.532
r209 106 107 1.86822 $w=3.87e-07 $l=1.5e-08 $layer=POLY_cond $X=3.425 $Y=1.532
+ $X2=3.44 $Y2=1.532
r210 104 105 7.83639 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.897 $Y=1.465
+ $X2=2.897 $Y2=1.63
r211 102 104 13.1437 $w=4.53e-07 $l=5e-07 $layer=LI1_cond $X=2.897 $Y=0.965
+ $X2=2.897 $Y2=1.465
r212 93 120 37.3643 $w=3.87e-07 $l=3e-07 $layer=POLY_cond $X=5.895 $Y=1.532
+ $X2=6.195 $Y2=1.532
r213 93 118 18.6822 $w=3.87e-07 $l=1.5e-07 $layer=POLY_cond $X=5.895 $Y=1.532
+ $X2=5.745 $Y2=1.532
r214 92 93 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=5.895
+ $Y=1.465 $X2=5.895 $Y2=1.465
r215 90 109 42.3463 $w=3.87e-07 $l=3.4e-07 $layer=POLY_cond $X=3.515 $Y=1.532
+ $X2=3.855 $Y2=1.532
r216 90 107 9.34109 $w=3.87e-07 $l=7.5e-08 $layer=POLY_cond $X=3.515 $Y=1.532
+ $X2=3.44 $Y2=1.532
r217 89 92 83.1156 $w=3.28e-07 $l=2.38e-06 $layer=LI1_cond $X=3.515 $Y=1.465
+ $X2=5.895 $Y2=1.465
r218 89 90 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=3.515
+ $Y=1.465 $X2=3.515 $Y2=1.465
r219 87 104 2.61955 $w=3.3e-07 $l=2.28e-07 $layer=LI1_cond $X=3.125 $Y=1.465
+ $X2=2.897 $Y2=1.465
r220 87 89 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.125 $Y=1.465
+ $X2=3.515 $Y2=1.465
r221 86 100 3.46198 $w=2.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=2.775 $Y=1.82
+ $X2=2.715 $Y2=1.905
r222 86 105 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=1.82
+ $X2=2.775 $Y2=1.63
r223 81 100 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=1.99
+ $X2=2.715 $Y2=1.905
r224 81 83 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=2.715 $Y=1.99
+ $X2=2.715 $Y2=2.815
r225 80 96 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=1.905
+ $X2=1.815 $Y2=1.905
r226 79 100 3.05049 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=1.905
+ $X2=2.715 $Y2=1.905
r227 79 80 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.55 $Y=1.905
+ $X2=1.98 $Y2=1.905
r228 78 98 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.935 $Y=1.005
+ $X2=1.81 $Y2=1.005
r229 78 102 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=1.935 $Y=1.005
+ $X2=2.67 $Y2=1.005
r230 73 98 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=0.88
+ $X2=1.81 $Y2=1.005
r231 73 75 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.81 $Y=0.88
+ $X2=1.81 $Y2=0.515
r232 69 96 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=1.99
+ $X2=1.815 $Y2=1.905
r233 69 71 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=1.815 $Y=1.99
+ $X2=1.815 $Y2=2.815
r234 66 123 25.0561 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.645 $Y=1.765
+ $X2=6.645 $Y2=1.532
r235 66 68 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.645 $Y=1.765
+ $X2=6.645 $Y2=2.4
r236 62 122 25.0561 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.635 $Y=1.3
+ $X2=6.635 $Y2=1.532
r237 62 64 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.635 $Y=1.3
+ $X2=6.635 $Y2=0.74
r238 58 121 25.0561 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.205 $Y=1.3
+ $X2=6.205 $Y2=1.532
r239 58 60 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.205 $Y=1.3
+ $X2=6.205 $Y2=0.74
r240 55 120 25.0561 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=1.532
r241 55 57 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=2.4
r242 52 118 25.0561 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=1.532
r243 52 54 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=2.4
r244 48 117 25.0561 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.705 $Y=1.3
+ $X2=5.705 $Y2=1.532
r245 48 50 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.705 $Y=1.3
+ $X2=5.705 $Y2=0.74
r246 45 116 25.0561 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.295 $Y=1.765
+ $X2=5.295 $Y2=1.532
r247 45 47 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.295 $Y=1.765
+ $X2=5.295 $Y2=2.4
r248 41 115 25.0561 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.215 $Y=1.3
+ $X2=5.215 $Y2=1.532
r249 41 43 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.215 $Y=1.3
+ $X2=5.215 $Y2=0.74
r250 38 114 25.0561 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.84 $Y=1.765
+ $X2=4.84 $Y2=1.532
r251 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.84 $Y=1.765
+ $X2=4.84 $Y2=2.4
r252 34 113 25.0561 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=1.532
r253 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=0.74
r254 31 112 25.0561 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.39 $Y=1.765
+ $X2=4.39 $Y2=1.532
r255 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.39 $Y=1.765
+ $X2=4.39 $Y2=2.4
r256 27 111 25.0561 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=1.532
r257 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=0.74
r258 24 110 25.0561 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.94 $Y=1.765
+ $X2=3.94 $Y2=1.532
r259 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.94 $Y=1.765
+ $X2=3.94 $Y2=2.4
r260 20 109 25.0561 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.855 $Y=1.3
+ $X2=3.855 $Y2=1.532
r261 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.855 $Y=1.3
+ $X2=3.855 $Y2=0.74
r262 17 107 25.0561 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.44 $Y=1.765
+ $X2=3.44 $Y2=1.532
r263 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.44 $Y=1.765
+ $X2=3.44 $Y2=2.4
r264 13 106 25.0561 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.425 $Y=1.3
+ $X2=3.425 $Y2=1.532
r265 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.425 $Y=1.3
+ $X2=3.425 $Y2=0.74
r266 4 100 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=1.84 $X2=2.715 $Y2=1.985
r267 4 83 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=1.84 $X2=2.715 $Y2=2.815
r268 3 96 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.84 $X2=1.815 $Y2=1.985
r269 3 71 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.84 $X2=1.815 $Y2=2.815
r270 2 102 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.37 $X2=2.71 $Y2=0.965
r271 1 98 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.37 $X2=1.85 $Y2=0.965
r272 1 75 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.37 $X2=1.85 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFBUF_8%VPWR 1 2 3 4 5 6 7 24 28 30 34 38 42 46 50
+ 52 54 58 60 65 70 75 80 86 89 92 95 98 101 105
r109 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r110 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r111 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r112 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r113 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 84 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r118 84 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r119 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r120 81 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.105 $Y=3.33
+ $X2=5.97 $Y2=3.33
r121 81 83 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.105 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 80 104 4.41691 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=6.967 $Y2=3.33
r123 80 83 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 79 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r125 79 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r126 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r127 76 98 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.067 $Y2=3.33
r128 76 78 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.52 $Y2=3.33
r129 75 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.97 $Y2=3.33
r130 75 78 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.52 $Y2=3.33
r131 74 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r132 74 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r134 71 95 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.162 $Y2=3.33
r135 71 73 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 70 98 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.93 $Y=3.33
+ $X2=5.067 $Y2=3.33
r137 70 73 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.93 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 69 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r139 69 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r141 66 86 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=0.742 $Y2=3.33
r142 66 68 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r143 65 89 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.265 $Y2=3.33
r144 65 68 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=1.2 $Y2=3.33
r145 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r146 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r147 60 86 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.742 $Y2=3.33
r148 60 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r149 58 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r150 58 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r151 54 57 26.4495 $w=3.03e-07 $l=7e-07 $layer=LI1_cond $X=6.887 $Y=2.115
+ $X2=6.887 $Y2=2.815
r152 52 104 3.14133 $w=3.05e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.887 $Y=3.245
+ $X2=6.967 $Y2=3.33
r153 52 57 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=6.887 $Y=3.245
+ $X2=6.887 $Y2=2.815
r154 48 101 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=3.245
+ $X2=5.97 $Y2=3.33
r155 48 50 40.1221 $w=2.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.97 $Y=3.245
+ $X2=5.97 $Y2=2.305
r156 44 98 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.067 $Y=3.245
+ $X2=5.067 $Y2=3.33
r157 44 46 39.3926 $w=2.73e-07 $l=9.4e-07 $layer=LI1_cond $X=5.067 $Y=3.245
+ $X2=5.067 $Y2=2.305
r158 40 95 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.162 $Y=3.245
+ $X2=4.162 $Y2=3.33
r159 40 42 42.4822 $w=2.53e-07 $l=9.4e-07 $layer=LI1_cond $X=4.162 $Y=3.245
+ $X2=4.162 $Y2=2.305
r160 39 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=3.33
+ $X2=3.215 $Y2=3.33
r161 38 95 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=4.162 $Y2=3.33
r162 38 39 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=3.38 $Y2=3.33
r163 34 37 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.215 $Y=1.985
+ $X2=3.215 $Y2=2.815
r164 32 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=3.245
+ $X2=3.215 $Y2=3.33
r165 32 37 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.215 $Y=3.245
+ $X2=3.215 $Y2=2.815
r166 31 89 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.265 $Y2=3.33
r167 30 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=3.215 $Y2=3.33
r168 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=2.38 $Y2=3.33
r169 26 89 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.265 $Y=3.245
+ $X2=2.265 $Y2=3.33
r170 26 28 46.0977 $w=2.28e-07 $l=9.2e-07 $layer=LI1_cond $X=2.265 $Y=3.245
+ $X2=2.265 $Y2=2.325
r171 22 86 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.742 $Y=3.245
+ $X2=0.742 $Y2=3.33
r172 22 24 23.0489 $w=3.53e-07 $l=7.1e-07 $layer=LI1_cond $X=0.742 $Y=3.245
+ $X2=0.742 $Y2=2.535
r173 7 57 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=6.72
+ $Y=1.84 $X2=6.875 $Y2=2.815
r174 7 54 400 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=6.72
+ $Y=1.84 $X2=6.875 $Y2=2.115
r175 6 50 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=5.82
+ $Y=1.84 $X2=5.97 $Y2=2.305
r176 5 46 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=4.915
+ $Y=1.84 $X2=5.065 $Y2=2.305
r177 4 42 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=4.015
+ $Y=1.84 $X2=4.165 $Y2=2.305
r178 3 37 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=1.84 $X2=3.215 $Y2=2.815
r179 3 34 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=1.84 $X2=3.215 $Y2=1.985
r180 2 28 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=2.115
+ $Y=1.84 $X2=2.265 $Y2=2.325
r181 1 24 600 $w=1.7e-07 $l=7.7086e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.74 $Y2=2.535
.ends

.subckt PM_SKY130_FD_SC_HS__BUFBUF_8%X 1 2 3 4 5 6 7 8 27 31 35 36 41 42 45 49
+ 53 57 61 63 65 69 70 71 75
r110 71 75 7.80543 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.96 $Y=1.665
+ $X2=6.665 $Y2=1.665
r111 65 67 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=6.42 $Y=1.985
+ $X2=6.42 $Y2=2.815
r112 63 65 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.42 $Y=1.97
+ $X2=6.42 $Y2=1.985
r113 59 61 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=6.42 $Y=0.88
+ $X2=6.42 $Y2=0.515
r114 58 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.655 $Y=1.885
+ $X2=5.52 $Y2=1.885
r115 57 63 5.08453 $w=5.54e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.255 $Y=1.885
+ $X2=6.42 $Y2=1.97
r116 57 75 4.84477 $w=5.54e-07 $l=5.08232e-07 $layer=LI1_cond $X=6.255 $Y=1.885
+ $X2=6.665 $Y2=1.665
r117 57 58 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.255 $Y=1.885
+ $X2=5.655 $Y2=1.885
r118 53 55 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=5.52 $Y=1.985
+ $X2=5.52 $Y2=2.815
r119 51 70 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=1.97
+ $X2=5.52 $Y2=1.885
r120 51 53 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.52 $Y=1.97
+ $X2=5.52 $Y2=1.985
r121 50 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.745 $Y=1.885
+ $X2=4.62 $Y2=1.885
r122 49 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.385 $Y=1.885
+ $X2=5.52 $Y2=1.885
r123 49 50 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.385 $Y=1.885
+ $X2=4.745 $Y2=1.885
r124 45 47 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.62 $Y=1.985
+ $X2=4.62 $Y2=2.815
r125 43 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=1.97
+ $X2=4.62 $Y2=1.885
r126 43 45 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=4.62 $Y=1.97
+ $X2=4.62 $Y2=1.985
r127 41 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.495 $Y=1.885
+ $X2=4.62 $Y2=1.885
r128 41 42 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.495 $Y=1.885
+ $X2=3.83 $Y2=1.885
r129 38 40 41.027 $w=2.48e-07 $l=8.9e-07 $layer=LI1_cond $X=4.57 $Y=1.005
+ $X2=5.46 $Y2=1.005
r130 36 38 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=3.805 $Y=1.005
+ $X2=4.57 $Y2=1.005
r131 35 75 14.5343 $w=5.54e-07 $l=8.40357e-07 $layer=LI1_cond $X=6.255 $Y=1.005
+ $X2=6.665 $Y2=1.665
r132 35 59 4.73129 $w=5.54e-07 $l=2.18746e-07 $layer=LI1_cond $X=6.255 $Y=1.005
+ $X2=6.42 $Y2=0.88
r133 35 40 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=6.255 $Y=1.005
+ $X2=5.46 $Y2=1.005
r134 31 33 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=3.697 $Y=1.985
+ $X2=3.697 $Y2=2.815
r135 29 42 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=3.697 $Y=1.97
+ $X2=3.83 $Y2=1.885
r136 29 31 0.652326 $w=2.63e-07 $l=1.5e-08 $layer=LI1_cond $X=3.697 $Y=1.97
+ $X2=3.697 $Y2=1.985
r137 25 36 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.64 $Y=0.88
+ $X2=3.805 $Y2=1.005
r138 25 27 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.64 $Y=0.88
+ $X2=3.64 $Y2=0.515
r139 8 67 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.84 $X2=6.42 $Y2=2.815
r140 8 65 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.84 $X2=6.42 $Y2=1.985
r141 7 55 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.37
+ $Y=1.84 $X2=5.52 $Y2=2.815
r142 7 53 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.37
+ $Y=1.84 $X2=5.52 $Y2=1.985
r143 6 47 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.465
+ $Y=1.84 $X2=4.615 $Y2=2.815
r144 6 45 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.465
+ $Y=1.84 $X2=4.615 $Y2=1.985
r145 5 33 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.84 $X2=3.715 $Y2=2.815
r146 5 31 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.84 $X2=3.715 $Y2=1.985
r147 4 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.28
+ $Y=0.37 $X2=6.42 $Y2=0.515
r148 3 40 182 $w=1.7e-07 $l=6.74667e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.37 $X2=5.46 $Y2=0.965
r149 2 38 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.965
r150 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.5
+ $Y=0.37 $X2=3.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFBUF_8%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48
+ 50 52 57 62 67 72 77 82 88 91 94 97 100 103 107
r101 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r102 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r103 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r104 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r105 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r106 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r107 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r108 86 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r109 86 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r110 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r111 83 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=0
+ $X2=5.92 $Y2=0
r112 83 85 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=0
+ $X2=6.48 $Y2=0
r113 82 106 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.977 $Y2=0
r114 82 85 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.48 $Y2=0
r115 81 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r116 81 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r117 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r118 78 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r119 78 80 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r120 77 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=5.92 $Y2=0
r121 77 80 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=5.52 $Y2=0
r122 76 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r123 76 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r124 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r125 73 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.14
+ $Y2=0
r126 73 75 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.305 $Y=0
+ $X2=4.56 $Y2=0
r127 72 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r128 72 75 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.56 $Y2=0
r129 68 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.14
+ $Y2=0
r130 68 70 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.6
+ $Y2=0
r131 67 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=4.14
+ $Y2=0
r132 67 70 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.6
+ $Y2=0
r133 66 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r134 66 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r135 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r136 63 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.28
+ $Y2=0
r137 63 65 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.64 $Y2=0
r138 62 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.14
+ $Y2=0
r139 62 65 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=2.64 $Y2=0
r140 61 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r141 61 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r142 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r143 58 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r144 58 60 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r145 57 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.28
+ $Y2=0
r146 57 60 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=1.2
+ $Y2=0
r147 55 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r148 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r149 52 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r150 52 54 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r151 50 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r152 50 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r153 50 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r154 46 106 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r155 46 48 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r156 42 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r157 42 44 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.545
r158 38 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r159 38 40 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.545
r160 34 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r161 34 36 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.545
r162 30 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r163 30 32 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.545
r164 26 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r165 26 28 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.545
r166 22 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r167 22 24 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.675
r168 7 48 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.71
+ $Y=0.37 $X2=6.92 $Y2=0.515
r169 6 44 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=5.78
+ $Y=0.37 $X2=5.92 $Y2=0.545
r170 5 40 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.545
r171 4 36 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.14 $Y2=0.545
r172 3 32 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.37 $X2=3.14 $Y2=0.545
r173 2 28 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.37 $X2=2.28 $Y2=0.545
r174 1 24 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.79 $Y2=0.675
.ends

