* File: sky130_fd_sc_hs__dlymetal6s2s_1.pex.spice
* Created: Thu Aug 27 20:43:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%A 3 5 7 8 12
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.39
+ $Y=1.44 $X2=0.39 $Y2=1.44
r31 8 12 5.98039 $w=4.48e-07 $l=2.25e-07 $layer=LI1_cond $X=0.33 $Y=1.665
+ $X2=0.33 $Y2=1.44
r32 5 11 64.5325 $w=2.97e-07 $l=3.66367e-07 $layer=POLY_cond $X=0.49 $Y=1.765
+ $X2=0.402 $Y2=1.44
r33 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.49 $Y=1.765 $X2=0.49
+ $Y2=2.05
r34 1 11 38.5662 $w=2.97e-07 $l=2.00237e-07 $layer=POLY_cond $X=0.48 $Y=1.275
+ $X2=0.402 $Y2=1.44
r35 1 3 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.48 $Y=1.275
+ $X2=0.48 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%A_28_138# 1 2 9 11 13 14 16 18 19 21
+ 28
c64 18 0 1.94125e-19 $X=0.81 $Y=1.605
r65 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.955
+ $Y=1.44 $X2=0.955 $Y2=1.44
r66 29 31 18.9224 $w=2.45e-07 $l=3.8e-07 $layer=LI1_cond $X=0.882 $Y=1.06
+ $X2=0.882 $Y2=1.44
r67 26 28 7.56208 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.08
+ $X2=0.43 $Y2=2.08
r68 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=0.247 $Y=0.865
+ $X2=0.247 $Y2=1.06
r69 18 31 9.37148 $w=2.45e-07 $l=1.9775e-07 $layer=LI1_cond $X=0.81 $Y=1.605
+ $X2=0.882 $Y2=1.44
r70 18 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.81 $Y=1.605
+ $X2=0.81 $Y2=1.935
r71 16 19 6.89401 $w=2.05e-07 $l=1.38109e-07 $layer=LI1_cond $X=0.725 $Y=2.037
+ $X2=0.81 $Y2=1.935
r72 16 28 15.9601 $w=2.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.725 $Y=2.037
+ $X2=0.43 $Y2=2.037
r73 15 23 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.395 $Y=1.06
+ $X2=0.247 $Y2=1.06
r74 14 29 2.87745 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=0.725 $Y=1.06
+ $X2=0.882 $Y2=1.06
r75 14 15 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.725 $Y=1.06
+ $X2=0.395 $Y2=1.06
r76 11 32 66.0502 $w=2.82e-07 $l=3.49106e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=0.955 $Y2=1.44
r77 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r78 7 32 41.2665 $w=2.82e-07 $l=1.8735e-07 $layer=POLY_cond $X=0.97 $Y=1.26
+ $X2=0.955 $Y2=1.44
r79 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.97 $Y=1.26 $X2=0.97
+ $Y2=0.74
r80 2 26 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.265 $Y2=2.06
r81 1 21 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.69 $X2=0.265 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%X 1 2 9 11 13 16 19 24 27 28 29 30 31
+ 37 39 45
c83 11 0 3.44873e-19 $X=1.975 $Y=1.765
r84 43 45 1.17953 $w=1.7e-07 $l=1.225e-06 $layer=MET1_cond $X=1.345 $Y=2.405
+ $X2=2.57 $Y2=2.405
r85 37 41 29.8172 $w=3.13e-07 $l=8.15e-07 $layer=LI1_cond $X=1.222 $Y=2
+ $X2=1.222 $Y2=2.815
r86 37 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035 $X2=1.2
+ $Y2=2.035
r87 31 43 0.0580243 $w=1.7e-07 $l=1.9e-07 $layer=MET1_cond $X=1.155 $Y=2.405
+ $X2=1.345 $Y2=2.405
r88 31 39 0.0820293 $w=7.6e-07 $l=2.85e-07 $layer=MET1_cond $X=1.155 $Y=2.32
+ $X2=1.155 $Y2=2.035
r89 31 45 0.199317 $w=1.7e-07 $l=2.07e-07 $layer=MET1_cond $X=2.777 $Y=2.405
+ $X2=2.57 $Y2=2.405
r90 27 37 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=1.222 $Y=1.992
+ $X2=1.222 $Y2=2
r91 27 28 8.16989 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=1.222 $Y=1.992
+ $X2=1.222 $Y2=1.835
r92 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.44 $X2=1.83 $Y2=1.44
r93 22 30 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=1.46
+ $X2=1.295 $Y2=1.46
r94 22 24 17.8827 $w=2.88e-07 $l=4.5e-07 $layer=LI1_cond $X=1.38 $Y=1.46
+ $X2=1.83 $Y2=1.46
r95 20 30 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.295 $Y=1.605
+ $X2=1.295 $Y2=1.46
r96 20 28 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.295 $Y=1.605
+ $X2=1.295 $Y2=1.835
r97 19 30 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.295 $Y=1.315
+ $X2=1.295 $Y2=1.46
r98 19 29 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.295 $Y=1.315
+ $X2=1.295 $Y2=1.075
r99 14 29 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.235 $Y=0.93
+ $X2=1.235 $Y2=1.075
r100 14 16 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=1.235 $Y=0.93
+ $X2=1.235 $Y2=0.57
r101 11 25 62.0998 $w=3.28e-07 $l=3.75999e-07 $layer=POLY_cond $X=1.975 $Y=1.765
+ $X2=1.865 $Y2=1.44
r102 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.975 $Y=1.765
+ $X2=1.975 $Y2=2.05
r103 7 25 38.5876 $w=3.28e-07 $l=1.90526e-07 $layer=POLY_cond $X=1.92 $Y=1.275
+ $X2=1.865 $Y2=1.44
r104 7 9 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.92 $Y=1.275
+ $X2=1.92 $Y2=0.9
r105 2 41 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=2.815
r106 2 37 400 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=2
r107 1 16 91 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.37 $X2=1.185 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%A_316_138# 1 2 9 11 13 14 16 18 19 21
+ 28
c65 11 0 3.02239e-19 $X=2.49 $Y=1.765
r66 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=1.44 $X2=2.44 $Y2=1.44
r67 26 28 4.97949 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.75 $Y=2.06
+ $X2=1.87 $Y2=2.06
r68 21 23 7.88514 $w=2.83e-07 $l=1.95e-07 $layer=LI1_cond $X=1.692 $Y=0.865
+ $X2=1.692 $Y2=1.06
r69 18 31 9.12826 $w=2.69e-07 $l=2.07123e-07 $layer=LI1_cond $X=2.25 $Y=1.605
+ $X2=2.345 $Y2=1.44
r70 18 19 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.25 $Y=1.605
+ $X2=2.25 $Y2=1.895
r71 16 19 7.11011 $w=2.45e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.165 $Y=2.017
+ $X2=2.25 $Y2=1.895
r72 16 28 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=2.165 $Y=2.017
+ $X2=1.87 $Y2=2.017
r73 15 23 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.835 $Y=1.06
+ $X2=1.692 $Y2=1.06
r74 14 31 17.2342 $w=2.69e-07 $l=4.61302e-07 $layer=LI1_cond $X=2.165 $Y=1.06
+ $X2=2.345 $Y2=1.44
r75 14 15 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.165 $Y=1.06
+ $X2=1.835 $Y2=1.06
r76 11 32 66.0502 $w=2.82e-07 $l=3.49106e-07 $layer=POLY_cond $X=2.49 $Y=1.765
+ $X2=2.44 $Y2=1.44
r77 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.49 $Y=1.765
+ $X2=2.49 $Y2=2.4
r78 7 32 41.2665 $w=2.82e-07 $l=1.94422e-07 $layer=POLY_cond $X=2.41 $Y=1.26
+ $X2=2.44 $Y2=1.44
r79 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.41 $Y=1.26 $X2=2.41
+ $Y2=0.74
r80 2 26 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=1.84 $X2=1.75 $Y2=2.06
r81 1 21 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.69 $X2=1.705 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%A_497_74# 1 2 9 11 13 16 20 23 28 31
+ 32 40 41
c65 40 0 1.50748e-19 $X=2.715 $Y=2
c66 11 0 1.53639e-19 $X=3.46 $Y=1.765
c67 9 0 1.48579e-19 $X=3.36 $Y=0.9
r68 40 42 5.47606 $w=3.58e-07 $l=1.6e-07 $layer=LI1_cond $X=2.685 $Y=2 $X2=2.685
+ $Y2=2.16
r69 40 41 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=2
+ $X2=2.685 $Y2=1.835
r70 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.44 $X2=3.27 $Y2=1.44
r71 26 32 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.46
+ $X2=2.78 $Y2=1.46
r72 26 28 16.0945 $w=2.88e-07 $l=4.05e-07 $layer=LI1_cond $X=2.865 $Y=1.46
+ $X2=3.27 $Y2=1.46
r73 24 32 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.78 $Y=1.605
+ $X2=2.78 $Y2=1.46
r74 24 41 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.78 $Y=1.605
+ $X2=2.78 $Y2=1.835
r75 23 32 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.78 $Y=1.315
+ $X2=2.78 $Y2=1.46
r76 23 31 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.78 $Y=1.315
+ $X2=2.78 $Y2=1.075
r77 20 42 25.1617 $w=2.98e-07 $l=6.55e-07 $layer=LI1_cond $X=2.715 $Y=2.815
+ $X2=2.715 $Y2=2.16
r78 14 31 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=2.697 $Y=0.908
+ $X2=2.697 $Y2=1.075
r79 14 16 11.6276 $w=3.33e-07 $l=3.38e-07 $layer=LI1_cond $X=2.697 $Y=0.908
+ $X2=2.697 $Y2=0.57
r80 11 29 60.4253 $w=3.58e-07 $l=3.85811e-07 $layer=POLY_cond $X=3.46 $Y=1.765
+ $X2=3.327 $Y2=1.44
r81 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.46 $Y=1.765
+ $X2=3.46 $Y2=2.05
r82 7 29 38.8834 $w=3.58e-07 $l=1.80748e-07 $layer=POLY_cond $X=3.36 $Y=1.275
+ $X2=3.327 $Y2=1.44
r83 7 9 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=3.36 $Y=1.275
+ $X2=3.36 $Y2=0.9
r84 2 40 400 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=1.84 $X2=2.715 $Y2=2
r85 2 20 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=1.84 $X2=2.715 $Y2=2.815
r86 1 16 91 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.37 $X2=2.625 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%A_604_138# 1 2 9 11 13 16 18 19 20 21
+ 23
r57 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.44 $X2=3.925 $Y2=1.44
r58 23 24 20.2615 $w=2.83e-07 $l=4.7e-07 $layer=LI1_cond $X=3.235 $Y=2.06
+ $X2=3.705 $Y2=2.06
r59 21 24 2.77065 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=1.895
+ $X2=3.705 $Y2=2.06
r60 20 27 8.10771 $w=2.93e-07 $l=2.09893e-07 $layer=LI1_cond $X=3.705 $Y=1.605
+ $X2=3.807 $Y2=1.44
r61 20 21 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=3.705 $Y=1.605
+ $X2=3.705 $Y2=1.895
r62 18 27 15.8225 $w=2.93e-07 $l=4.70277e-07 $layer=LI1_cond $X=3.605 $Y=1.06
+ $X2=3.807 $Y2=1.44
r63 18 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.605 $Y=1.06
+ $X2=3.275 $Y2=1.06
r64 14 19 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=3.167 $Y=0.975
+ $X2=3.275 $Y2=1.06
r65 14 16 5.89622 $w=2.13e-07 $l=1.1e-07 $layer=LI1_cond $X=3.167 $Y=0.975
+ $X2=3.167 $Y2=0.865
r66 11 28 66.0502 $w=2.82e-07 $l=3.51426e-07 $layer=POLY_cond $X=3.98 $Y=1.765
+ $X2=3.925 $Y2=1.44
r67 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.98 $Y=1.765
+ $X2=3.98 $Y2=2.4
r68 7 28 41.2665 $w=2.82e-07 $l=2.14243e-07 $layer=POLY_cond $X=3.85 $Y=1.26
+ $X2=3.925 $Y2=1.44
r69 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.85 $Y=1.26 $X2=3.85
+ $Y2=0.74
r70 2 23 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=1.84 $X2=3.235 $Y2=2.06
r71 1 16 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.69 $X2=3.145 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%VPWR 1 2 3 12 16 20 22 24 29 34 41 42
+ 45 48 51 58
r50 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r51 49 58 0.0655027 $w=4.9e-07 $l=2.35e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.925 $Y2=3.33
r52 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 42 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 39 51 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=3.732 $Y2=3.33
r57 39 41 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 38 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 35 48 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.247 $Y2=3.33
r61 35 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 34 51 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=3.732 $Y2=3.33
r63 34 37 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 33 58 0.202083 $w=4.9e-07 $l=7.25e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.925 $Y2=3.33
r65 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r67 30 45 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.737 $Y2=3.33
r68 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 29 48 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.1 $Y=3.33
+ $X2=2.247 $Y2=3.33
r70 29 32 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.1 $Y=3.33 $X2=1.2
+ $Y2=3.33
r71 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r73 24 45 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.737 $Y2=3.33
r74 24 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.24 $Y2=3.33
r75 22 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r76 22 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 18 51 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.732 $Y=3.245
+ $X2=3.732 $Y2=3.33
r78 18 20 30.0807 $w=2.93e-07 $l=7.7e-07 $layer=LI1_cond $X=3.732 $Y=3.245
+ $X2=3.732 $Y2=2.475
r79 14 48 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.247 $Y=3.245
+ $X2=2.247 $Y2=3.33
r80 14 16 30.0807 $w=2.93e-07 $l=7.7e-07 $layer=LI1_cond $X=2.247 $Y=3.245
+ $X2=2.247 $Y2=2.475
r81 10 45 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.737 $Y=3.245
+ $X2=0.737 $Y2=3.33
r82 10 12 30.0807 $w=2.93e-07 $l=7.7e-07 $layer=LI1_cond $X=0.737 $Y=3.245
+ $X2=0.737 $Y2=2.475
r83 3 20 300 $w=1.7e-07 $l=7.34677e-07 $layer=licon1_PDIFF $count=2 $X=3.535
+ $Y=1.84 $X2=3.75 $Y2=2.475
r84 2 16 300 $w=1.7e-07 $l=7.34677e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=1.84 $X2=2.265 $Y2=2.475
r85 1 12 300 $w=1.7e-07 $l=7.34677e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.84 $X2=0.78 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%A_785_74# 1 2 9 13 17 24 25
c31 24 0 1.53639e-19 $X=4.205 $Y=2
r32 24 26 5.41124 $w=3.73e-07 $l=1.6e-07 $layer=LI1_cond $X=4.162 $Y=2 $X2=4.162
+ $Y2=2.16
r33 24 25 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=4.162 $Y=2
+ $X2=4.162 $Y2=1.835
r34 17 25 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.265 $Y=1.075
+ $X2=4.265 $Y2=1.835
r35 13 26 25.1617 $w=2.98e-07 $l=6.55e-07 $layer=LI1_cond $X=4.2 $Y=2.815
+ $X2=4.2 $Y2=2.16
r36 7 17 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=4.16 $Y=0.885
+ $X2=4.16 $Y2=1.075
r37 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=4.16 $Y=0.885
+ $X2=4.16 $Y2=0.57
r38 2 24 400 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.84 $X2=4.205 $Y2=2
r39 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.84 $X2=4.205 $Y2=2.815
r40 1 9 91 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=2 $X=3.925
+ $Y=0.37 $X2=4.065 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__DLYMETAL6S2S_1%VGND 1 2 3 12 16 20 22 24 29 34 41 42
+ 45 48 51 58
c59 16 0 1.5366e-19 $X=2.195 $Y=0.72
r60 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r61 49 58 0.0655027 $w=4.9e-07 $l=2.35e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.925 $Y2=0
r62 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r64 42 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r65 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=3.635
+ $Y2=0
r67 39 41 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=4.56
+ $Y2=0
r68 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r69 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r70 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.195
+ $Y2=0
r71 35 37 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=3.12
+ $Y2=0
r72 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.635
+ $Y2=0
r73 34 37 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.12
+ $Y2=0
r74 33 58 0.06829 $w=4.9e-07 $l=2.45e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.925
+ $Y2=0
r75 33 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r76 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r77 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=0.755
+ $Y2=0
r78 30 32 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=1.68
+ $Y2=0
r79 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.195
+ $Y2=0
r80 29 32 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.68
+ $Y2=0
r81 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r82 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r83 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.755
+ $Y2=0
r84 24 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.24
+ $Y2=0
r85 22 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r86 22 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r87 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0.085
+ $X2=3.635 $Y2=0
r88 18 20 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.635 $Y=0.085
+ $X2=3.635 $Y2=0.72
r89 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0
r90 14 16 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0.72
r91 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r92 10 12 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.72
r93 3 20 182 $w=1.7e-07 $l=2.14476e-07 $layer=licon1_NDIFF $count=1 $X=3.435
+ $Y=0.69 $X2=3.635 $Y2=0.72
r94 2 16 182 $w=1.7e-07 $l=2.14476e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.69 $X2=2.195 $Y2=0.72
r95 1 12 182 $w=1.7e-07 $l=2.14476e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.69 $X2=0.755 $Y2=0.72
.ends

