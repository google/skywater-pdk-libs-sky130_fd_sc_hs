* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__fah_2 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_481_379# B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.948e+11p pd=2.99e+06u as=2.5648e+12p ps=2.029e+07u
M1001 a_1689_424# CI VPWR VPB pshort w=1e+06u l=150000u
+  ad=1.0242e+12p pd=6.01e+06u as=0p ps=0u
M1002 a_114_368# a_81_260# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=7e+11p pd=5.4e+06u as=0p ps=0u
M1003 a_514_424# a_481_379# a_413_392# VPB pshort w=840000u l=150000u
+  ad=7.686e+11p pd=3.51e+06u as=5.8e+11p ps=4.96e+06u
M1004 a_1689_424# a_849_424# a_1451_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=8.736e+11p ps=3.76e+06u
M1005 a_413_392# A VGND VNB nlowvt w=640000u l=150000u
+  ad=4.247e+11p pd=4.22e+06u as=1.82425e+12p ps=1.593e+07u
M1006 a_514_424# B a_413_392# VNB nlowvt w=640000u l=150000u
+  ad=3.904e+11p pd=2.5e+06u as=0p ps=0u
M1007 a_849_424# B a_114_368# VNB nlowvt w=640000u l=150000u
+  ad=4.448e+11p pd=2.67e+06u as=7.401e+11p ps=4.99e+06u
M1008 a_114_368# a_481_379# a_514_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1895_424# a_849_424# a_1689_424# VNB nlowvt w=640000u l=150000u
+  ad=4.729e+11p pd=2.9e+06u as=6.112e+11p ps=4.47e+06u
M1010 a_114_368# B a_514_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_1689_424# a_2052_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.12e+06u
M1012 a_1451_424# a_514_424# a_481_379# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_2052_424# a_849_424# a_1895_424# VPB pshort w=840000u l=150000u
+  ad=4.918e+11p pd=3.07e+06u as=5.334e+11p ps=2.95e+06u
M1014 COUT a_1451_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1015 VPWR A a_81_260# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1016 a_849_424# a_481_379# a_114_368# VPB pshort w=840000u l=150000u
+  ad=1.1298e+12p pd=4.37e+06u as=0p ps=0u
M1017 VGND A a_81_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.272e+11p ps=1.99e+06u
M1018 VPWR a_1895_424# SUM VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.472e+11p ps=2.86e+06u
M1019 a_1451_424# a_849_424# a_481_379# VNB nlowvt w=640000u l=150000u
+  ad=5.6e+11p pd=3.03e+06u as=2.33e+11p ps=2.13e+06u
M1020 a_1689_424# a_514_424# a_1451_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1689_424# CI VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1895_424# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.146e+11p ps=2.06e+06u
M1023 COUT a_1451_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1024 a_413_392# B a_849_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_413_392# a_481_379# a_849_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1451_424# COUT VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_2052_424# a_514_424# a_1895_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 SUM a_1895_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 SUM a_1895_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_413_392# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1895_424# a_514_424# a_1689_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_1689_424# a_2052_424# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_481_379# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_114_368# a_81_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_1451_424# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
